module day05_checker (
    valid,
    clear,
    clock,
    ingredient_id,
    is_fresh,
    total_count
);

    input valid;
    input clear;
    input clock;
    input [63:0] ingredient_id;
    output is_fresh;
    output [63:0] total_count;

    wire _2;
    wire _1697;
    wire [63:0] _13;
    wire _4;
    wire _6;
    wire [63:0] _1699;
    wire [63:0] _1700;
    wire [63:0] _7;
    reg [63:0] _1698;
    wire [64:0] _1692;
    wire _1693;
    wire _1694;
    wire [64:0] _1689;
    wire [64:0] _1688;
    wire _1690;
    wire _1691;
    wire _1695;
    wire [64:0] _1683;
    wire _1684;
    wire _1685;
    wire [64:0] _1680;
    wire [64:0] _1679;
    wire _1681;
    wire _1682;
    wire _1686;
    wire [64:0] _1674;
    wire _1675;
    wire _1676;
    wire [64:0] _1671;
    wire [64:0] _1670;
    wire _1672;
    wire _1673;
    wire _1677;
    wire [64:0] _1665;
    wire _1666;
    wire _1667;
    wire [64:0] _1662;
    wire [64:0] _1661;
    wire _1663;
    wire _1664;
    wire _1668;
    wire [64:0] _1656;
    wire _1657;
    wire _1658;
    wire [64:0] _1653;
    wire [64:0] _1652;
    wire _1654;
    wire _1655;
    wire _1659;
    wire [64:0] _1647;
    wire _1648;
    wire _1649;
    wire [64:0] _1644;
    wire [64:0] _1643;
    wire _1645;
    wire _1646;
    wire _1650;
    wire [64:0] _1638;
    wire _1639;
    wire _1640;
    wire [64:0] _1635;
    wire [64:0] _1634;
    wire _1636;
    wire _1637;
    wire _1641;
    wire [64:0] _1629;
    wire _1630;
    wire _1631;
    wire [64:0] _1626;
    wire [64:0] _1625;
    wire _1627;
    wire _1628;
    wire _1632;
    wire [64:0] _1620;
    wire _1621;
    wire _1622;
    wire [64:0] _1617;
    wire [64:0] _1616;
    wire _1618;
    wire _1619;
    wire _1623;
    wire [64:0] _1611;
    wire _1612;
    wire _1613;
    wire [64:0] _1608;
    wire [64:0] _1607;
    wire _1609;
    wire _1610;
    wire _1614;
    wire [64:0] _1602;
    wire _1603;
    wire _1604;
    wire [64:0] _1599;
    wire [64:0] _1598;
    wire _1600;
    wire _1601;
    wire _1605;
    wire [64:0] _1593;
    wire _1594;
    wire _1595;
    wire [64:0] _1590;
    wire [64:0] _1589;
    wire _1591;
    wire _1592;
    wire _1596;
    wire [64:0] _1584;
    wire _1585;
    wire _1586;
    wire [64:0] _1581;
    wire [64:0] _1580;
    wire _1582;
    wire _1583;
    wire _1587;
    wire [64:0] _1575;
    wire _1576;
    wire _1577;
    wire [64:0] _1572;
    wire [64:0] _1571;
    wire _1573;
    wire _1574;
    wire _1578;
    wire [64:0] _1566;
    wire _1567;
    wire _1568;
    wire [64:0] _1562;
    wire _1564;
    wire _1565;
    wire _1569;
    wire [64:0] _1557;
    wire _1558;
    wire _1559;
    wire [64:0] _1554;
    wire [64:0] _1553;
    wire _1555;
    wire _1556;
    wire _1560;
    wire [64:0] _1548;
    wire _1549;
    wire _1550;
    wire [64:0] _1545;
    wire [64:0] _1544;
    wire _1546;
    wire _1547;
    wire _1551;
    wire [64:0] _1539;
    wire _1540;
    wire _1541;
    wire [64:0] _1536;
    wire [64:0] _1535;
    wire _1537;
    wire _1538;
    wire _1542;
    wire [64:0] _1530;
    wire _1531;
    wire _1532;
    wire [64:0] _1527;
    wire [64:0] _1526;
    wire _1528;
    wire _1529;
    wire _1533;
    wire [64:0] _1521;
    wire _1522;
    wire _1523;
    wire [64:0] _1517;
    wire _1519;
    wire _1520;
    wire _1524;
    wire [64:0] _1512;
    wire _1513;
    wire _1514;
    wire [64:0] _1509;
    wire [64:0] _1508;
    wire _1510;
    wire _1511;
    wire _1515;
    wire [64:0] _1503;
    wire _1504;
    wire _1505;
    wire [64:0] _1500;
    wire [64:0] _1499;
    wire _1501;
    wire _1502;
    wire _1506;
    wire [64:0] _1494;
    wire _1495;
    wire _1496;
    wire [64:0] _1491;
    wire [64:0] _1490;
    wire _1492;
    wire _1493;
    wire _1497;
    wire [64:0] _1485;
    wire _1486;
    wire _1487;
    wire [64:0] _1482;
    wire [64:0] _1481;
    wire _1483;
    wire _1484;
    wire _1488;
    wire [64:0] _1476;
    wire _1477;
    wire _1478;
    wire [64:0] _1473;
    wire [64:0] _1472;
    wire _1474;
    wire _1475;
    wire _1479;
    wire [64:0] _1467;
    wire _1468;
    wire _1469;
    wire [64:0] _1464;
    wire [64:0] _1463;
    wire _1465;
    wire _1466;
    wire _1470;
    wire [64:0] _1458;
    wire _1459;
    wire _1460;
    wire [64:0] _1455;
    wire [64:0] _1454;
    wire _1456;
    wire _1457;
    wire _1461;
    wire [64:0] _1449;
    wire _1450;
    wire _1451;
    wire [64:0] _1446;
    wire [64:0] _1445;
    wire _1447;
    wire _1448;
    wire _1452;
    wire [64:0] _1440;
    wire _1441;
    wire _1442;
    wire [64:0] _1437;
    wire [64:0] _1436;
    wire _1438;
    wire _1439;
    wire _1443;
    wire [64:0] _1431;
    wire _1432;
    wire _1433;
    wire [64:0] _1428;
    wire [64:0] _1427;
    wire _1429;
    wire _1430;
    wire _1434;
    wire _1423;
    wire _1424;
    wire [64:0] _1419;
    wire [64:0] _1418;
    wire _1420;
    wire _1421;
    wire _1425;
    wire [64:0] _1413;
    wire _1414;
    wire _1415;
    wire [64:0] _1409;
    wire _1411;
    wire _1412;
    wire _1416;
    wire [64:0] _1404;
    wire _1405;
    wire _1406;
    wire [64:0] _1401;
    wire [64:0] _1400;
    wire _1402;
    wire _1403;
    wire _1407;
    wire [64:0] _1395;
    wire _1396;
    wire _1397;
    wire [64:0] _1391;
    wire _1393;
    wire _1394;
    wire _1398;
    wire [64:0] _1386;
    wire _1387;
    wire _1388;
    wire [64:0] _1383;
    wire [64:0] _1382;
    wire _1384;
    wire _1385;
    wire _1389;
    wire [64:0] _1377;
    wire _1378;
    wire _1379;
    wire [64:0] _1374;
    wire [64:0] _1373;
    wire _1375;
    wire _1376;
    wire _1380;
    wire [64:0] _1368;
    wire _1369;
    wire _1370;
    wire [64:0] _1365;
    wire [64:0] _1364;
    wire _1366;
    wire _1367;
    wire _1371;
    wire [64:0] _1359;
    wire _1360;
    wire _1361;
    wire [64:0] _1356;
    wire [64:0] _1355;
    wire _1357;
    wire _1358;
    wire _1362;
    wire [64:0] _1350;
    wire _1351;
    wire _1352;
    wire [64:0] _1347;
    wire [64:0] _1346;
    wire _1348;
    wire _1349;
    wire _1353;
    wire [64:0] _1341;
    wire _1342;
    wire _1343;
    wire [64:0] _1337;
    wire _1339;
    wire _1340;
    wire _1344;
    wire [64:0] _1332;
    wire _1333;
    wire _1334;
    wire [64:0] _1329;
    wire [64:0] _1328;
    wire _1330;
    wire _1331;
    wire _1335;
    wire [64:0] _1323;
    wire _1324;
    wire _1325;
    wire [64:0] _1320;
    wire [64:0] _1319;
    wire _1321;
    wire _1322;
    wire _1326;
    wire [64:0] _1314;
    wire _1315;
    wire _1316;
    wire [64:0] _1311;
    wire [64:0] _1310;
    wire _1312;
    wire _1313;
    wire _1317;
    wire [64:0] _1305;
    wire _1306;
    wire _1307;
    wire [64:0] _1302;
    wire [64:0] _1301;
    wire _1303;
    wire _1304;
    wire _1308;
    wire _1297;
    wire _1298;
    wire [64:0] _1293;
    wire [64:0] _1292;
    wire _1294;
    wire _1295;
    wire _1299;
    wire [64:0] _1287;
    wire _1288;
    wire _1289;
    wire [64:0] _1283;
    wire _1285;
    wire _1286;
    wire _1290;
    wire [64:0] _1278;
    wire _1279;
    wire _1280;
    wire [64:0] _1275;
    wire [64:0] _1274;
    wire _1276;
    wire _1277;
    wire _1281;
    wire [64:0] _1269;
    wire _1270;
    wire _1271;
    wire [64:0] _1265;
    wire _1267;
    wire _1268;
    wire _1272;
    wire [64:0] _1260;
    wire _1261;
    wire _1262;
    wire [64:0] _1256;
    wire _1258;
    wire _1259;
    wire _1263;
    wire [64:0] _1251;
    wire _1252;
    wire _1253;
    wire [64:0] _1248;
    wire [64:0] _1247;
    wire _1249;
    wire _1250;
    wire _1254;
    wire [64:0] _1242;
    wire _1243;
    wire _1244;
    wire [64:0] _1239;
    wire [64:0] _1238;
    wire _1240;
    wire _1241;
    wire _1245;
    wire [64:0] _1233;
    wire _1234;
    wire _1235;
    wire [64:0] _1230;
    wire [64:0] _1229;
    wire _1231;
    wire _1232;
    wire _1236;
    wire [64:0] _1224;
    wire _1225;
    wire _1226;
    wire [64:0] _1221;
    wire [64:0] _1220;
    wire _1222;
    wire _1223;
    wire _1227;
    wire [64:0] _1215;
    wire _1216;
    wire _1217;
    wire [64:0] _1212;
    wire [64:0] _1211;
    wire _1213;
    wire _1214;
    wire _1218;
    wire [64:0] _1206;
    wire _1207;
    wire _1208;
    wire [64:0] _1203;
    wire [64:0] _1202;
    wire _1204;
    wire _1205;
    wire _1209;
    wire _1198;
    wire _1199;
    wire [64:0] _1193;
    wire _1195;
    wire _1196;
    wire _1200;
    wire [64:0] _1188;
    wire _1189;
    wire _1190;
    wire [64:0] _1185;
    wire [64:0] _1184;
    wire _1186;
    wire _1187;
    wire _1191;
    wire [64:0] _1179;
    wire _1180;
    wire _1181;
    wire [64:0] _1175;
    wire _1177;
    wire _1178;
    wire _1182;
    wire [64:0] _1170;
    wire _1171;
    wire _1172;
    wire [64:0] _1167;
    wire [64:0] _1166;
    wire _1168;
    wire _1169;
    wire _1173;
    wire [64:0] _1161;
    wire _1162;
    wire _1163;
    wire [64:0] _1158;
    wire [64:0] _1157;
    wire _1159;
    wire _1160;
    wire _1164;
    wire [64:0] _1152;
    wire _1153;
    wire _1154;
    wire [64:0] _1149;
    wire [64:0] _1148;
    wire _1150;
    wire _1151;
    wire _1155;
    wire [64:0] _1143;
    wire _1144;
    wire _1145;
    wire [64:0] _1140;
    wire [64:0] _1139;
    wire _1141;
    wire _1142;
    wire _1146;
    wire [64:0] _1134;
    wire _1135;
    wire _1136;
    wire [64:0] _1131;
    wire [64:0] _1130;
    wire _1132;
    wire _1133;
    wire _1137;
    wire [64:0] _1125;
    wire _1126;
    wire _1127;
    wire [64:0] _1122;
    wire [64:0] _1121;
    wire _1123;
    wire _1124;
    wire _1128;
    wire [64:0] _1116;
    wire _1117;
    wire _1118;
    wire [64:0] _1113;
    wire [64:0] _1112;
    wire _1114;
    wire _1115;
    wire _1119;
    wire [64:0] _1107;
    wire _1108;
    wire _1109;
    wire [64:0] _1104;
    wire [64:0] _1103;
    wire _1105;
    wire _1106;
    wire _1110;
    wire [64:0] _1098;
    wire _1099;
    wire _1100;
    wire [64:0] _1095;
    wire [64:0] _1094;
    wire _1096;
    wire _1097;
    wire _1101;
    wire [64:0] _1089;
    wire _1090;
    wire _1091;
    wire [64:0] _1086;
    wire [64:0] _1085;
    wire _1087;
    wire _1088;
    wire _1092;
    wire [64:0] _1080;
    wire _1081;
    wire _1082;
    wire [64:0] _1077;
    wire [64:0] _1076;
    wire _1078;
    wire _1079;
    wire _1083;
    wire [64:0] _1071;
    wire _1072;
    wire _1073;
    wire [64:0] _1068;
    wire [64:0] _1067;
    wire _1069;
    wire _1070;
    wire _1074;
    wire [64:0] _1062;
    wire _1063;
    wire _1064;
    wire [64:0] _1059;
    wire [64:0] _1058;
    wire _1060;
    wire _1061;
    wire _1065;
    wire _1054;
    wire _1055;
    wire [64:0] _1049;
    wire _1051;
    wire _1052;
    wire _1056;
    wire [64:0] _1044;
    wire _1045;
    wire _1046;
    wire [64:0] _1041;
    wire [64:0] _1040;
    wire _1042;
    wire _1043;
    wire _1047;
    wire [64:0] _1035;
    wire _1036;
    wire _1037;
    wire [64:0] _1032;
    wire [64:0] _1031;
    wire _1033;
    wire _1034;
    wire _1038;
    wire [64:0] _1026;
    wire _1027;
    wire _1028;
    wire [64:0] _1023;
    wire [64:0] _1022;
    wire _1024;
    wire _1025;
    wire _1029;
    wire _1018;
    wire _1019;
    wire [64:0] _1014;
    wire [64:0] _1013;
    wire _1015;
    wire _1016;
    wire _1020;
    wire [64:0] _1008;
    wire _1009;
    wire _1010;
    wire [64:0] _1005;
    wire [64:0] _1004;
    wire _1006;
    wire _1007;
    wire _1011;
    wire [64:0] _999;
    wire _1000;
    wire _1001;
    wire [64:0] _996;
    wire [64:0] _995;
    wire _997;
    wire _998;
    wire _1002;
    wire [64:0] _990;
    wire _991;
    wire _992;
    wire [64:0] _986;
    wire _988;
    wire _989;
    wire _993;
    wire [64:0] _981;
    wire _982;
    wire _983;
    wire [64:0] _978;
    wire [64:0] _977;
    wire _979;
    wire _980;
    wire _984;
    wire [64:0] _972;
    wire _973;
    wire _974;
    wire [64:0] _969;
    wire [64:0] _968;
    wire _970;
    wire _971;
    wire _975;
    wire [64:0] _963;
    wire _964;
    wire _965;
    wire [64:0] _960;
    wire [64:0] _959;
    wire _961;
    wire _962;
    wire _966;
    wire [64:0] _954;
    wire _955;
    wire _956;
    wire [64:0] _951;
    wire [64:0] _950;
    wire _952;
    wire _953;
    wire _957;
    wire [64:0] _945;
    wire _946;
    wire _947;
    wire [64:0] _941;
    wire _943;
    wire _944;
    wire _948;
    wire [64:0] _936;
    wire _937;
    wire _938;
    wire [64:0] _933;
    wire [64:0] _932;
    wire _934;
    wire _935;
    wire _939;
    wire [64:0] _927;
    wire _928;
    wire _929;
    wire [64:0] _924;
    wire [64:0] _923;
    wire _925;
    wire _926;
    wire _930;
    wire [64:0] _918;
    wire _919;
    wire _920;
    wire [64:0] _914;
    wire _916;
    wire _917;
    wire _921;
    wire [64:0] _909;
    wire _910;
    wire _911;
    wire [64:0] _906;
    wire [64:0] _905;
    wire _907;
    wire _908;
    wire _912;
    wire [64:0] _900;
    wire _901;
    wire _902;
    wire [64:0] _897;
    wire [64:0] _896;
    wire _898;
    wire _899;
    wire _903;
    wire [64:0] _891;
    wire _892;
    wire _893;
    wire [64:0] _888;
    wire [64:0] _887;
    wire _889;
    wire _890;
    wire _894;
    wire [64:0] _882;
    wire _883;
    wire _884;
    wire [64:0] _879;
    wire [64:0] _878;
    wire _880;
    wire _881;
    wire _885;
    wire [64:0] _873;
    wire _874;
    wire _875;
    wire [64:0] _870;
    wire [64:0] _869;
    wire _871;
    wire _872;
    wire _876;
    wire [64:0] _864;
    wire _865;
    wire _866;
    wire [64:0] _861;
    wire [64:0] _860;
    wire _862;
    wire _863;
    wire _867;
    wire _856;
    wire _857;
    wire [64:0] _852;
    wire [64:0] _851;
    wire _853;
    wire _854;
    wire _858;
    wire [64:0] _846;
    wire _847;
    wire _848;
    wire [64:0] _843;
    wire [64:0] _842;
    wire _844;
    wire _845;
    wire _849;
    wire [64:0] _837;
    wire _838;
    wire _839;
    wire [64:0] _833;
    wire _835;
    wire _836;
    wire _840;
    wire _829;
    wire _830;
    wire [64:0] _824;
    wire _826;
    wire _827;
    wire _831;
    wire [64:0] _819;
    wire _820;
    wire _821;
    wire [64:0] _816;
    wire [64:0] _815;
    wire _817;
    wire _818;
    wire _822;
    wire [64:0] _810;
    wire _811;
    wire _812;
    wire [64:0] _807;
    wire [64:0] _806;
    wire _808;
    wire _809;
    wire _813;
    wire [64:0] _801;
    wire _802;
    wire _803;
    wire [64:0] _798;
    wire [64:0] _797;
    wire _799;
    wire _800;
    wire _804;
    wire [64:0] _792;
    wire _793;
    wire _794;
    wire [64:0] _789;
    wire [64:0] _788;
    wire _790;
    wire _791;
    wire _795;
    wire _784;
    wire _785;
    wire [64:0] _780;
    wire [64:0] _779;
    wire _781;
    wire _782;
    wire _786;
    wire [64:0] _774;
    wire _775;
    wire _776;
    wire [64:0] _771;
    wire [64:0] _770;
    wire _772;
    wire _773;
    wire _777;
    wire _766;
    wire _767;
    wire [64:0] _762;
    wire [64:0] _761;
    wire _763;
    wire _764;
    wire _768;
    wire [64:0] _756;
    wire _757;
    wire _758;
    wire [64:0] _753;
    wire [64:0] _752;
    wire _754;
    wire _755;
    wire _759;
    wire [64:0] _747;
    wire _748;
    wire _749;
    wire [64:0] _744;
    wire [64:0] _743;
    wire _745;
    wire _746;
    wire _750;
    wire [64:0] _738;
    wire _739;
    wire _740;
    wire [64:0] _735;
    wire [64:0] _734;
    wire _736;
    wire _737;
    wire _741;
    wire [64:0] _729;
    wire _730;
    wire _731;
    wire [64:0] _725;
    wire _727;
    wire _728;
    wire _732;
    wire [64:0] _720;
    wire _721;
    wire _722;
    wire [64:0] _717;
    wire [64:0] _716;
    wire _718;
    wire _719;
    wire _723;
    wire [64:0] _711;
    wire _712;
    wire _713;
    wire [64:0] _708;
    wire [64:0] _707;
    wire _709;
    wire _710;
    wire _714;
    wire [64:0] _702;
    wire _703;
    wire _704;
    wire [64:0] _698;
    wire _700;
    wire _701;
    wire _705;
    wire [64:0] _693;
    wire _694;
    wire _695;
    wire [64:0] _690;
    wire [64:0] _689;
    wire _691;
    wire _692;
    wire _696;
    wire [64:0] _684;
    wire _685;
    wire _686;
    wire [64:0] _681;
    wire [64:0] _680;
    wire _682;
    wire _683;
    wire _687;
    wire [64:0] _675;
    wire _676;
    wire _677;
    wire [64:0] _672;
    wire [64:0] _671;
    wire _673;
    wire _674;
    wire _678;
    wire [64:0] _666;
    wire _667;
    wire _668;
    wire [64:0] _662;
    wire _664;
    wire _665;
    wire _669;
    wire [64:0] _657;
    wire _658;
    wire _659;
    wire [64:0] _653;
    wire _655;
    wire _656;
    wire _660;
    wire [64:0] _648;
    wire _649;
    wire _650;
    wire [64:0] _645;
    wire [64:0] _644;
    wire _646;
    wire _647;
    wire _651;
    wire [64:0] _639;
    wire _640;
    wire _641;
    wire [64:0] _636;
    wire [64:0] _635;
    wire _637;
    wire _638;
    wire _642;
    wire [64:0] _630;
    wire _631;
    wire _632;
    wire [64:0] _626;
    wire _628;
    wire _629;
    wire _633;
    wire [64:0] _621;
    wire _622;
    wire _623;
    wire [64:0] _618;
    wire [64:0] _617;
    wire _619;
    wire _620;
    wire _624;
    wire [64:0] _612;
    wire _613;
    wire _614;
    wire [64:0] _609;
    wire [64:0] _608;
    wire _610;
    wire _611;
    wire _615;
    wire _604;
    wire _605;
    wire [64:0] _599;
    wire _601;
    wire _602;
    wire _606;
    wire _595;
    wire _596;
    wire [64:0] _591;
    wire [64:0] _590;
    wire _592;
    wire _593;
    wire _597;
    wire [64:0] _585;
    wire _586;
    wire _587;
    wire [64:0] _582;
    wire [64:0] _581;
    wire _583;
    wire _584;
    wire _588;
    wire [64:0] _576;
    wire _577;
    wire _578;
    wire [64:0] _573;
    wire [64:0] _572;
    wire _574;
    wire _575;
    wire _579;
    wire [64:0] _567;
    wire _568;
    wire _569;
    wire [64:0] _564;
    wire [64:0] _563;
    wire _565;
    wire _566;
    wire _570;
    wire _559;
    wire _560;
    wire [64:0] _554;
    wire _556;
    wire _557;
    wire _561;
    wire [64:0] _549;
    wire _550;
    wire _551;
    wire [64:0] _546;
    wire [64:0] _545;
    wire _547;
    wire _548;
    wire _552;
    wire _541;
    wire _542;
    wire [64:0] _536;
    wire _538;
    wire _539;
    wire _543;
    wire _532;
    wire _533;
    wire [64:0] _528;
    wire [64:0] _527;
    wire _529;
    wire _530;
    wire _534;
    wire [64:0] _522;
    wire _523;
    wire _524;
    wire [64:0] _519;
    wire [64:0] _518;
    wire _520;
    wire _521;
    wire _525;
    wire [64:0] _513;
    wire _514;
    wire _515;
    wire [64:0] _510;
    wire [64:0] _509;
    wire _511;
    wire _512;
    wire _516;
    wire _505;
    wire _506;
    wire [64:0] _500;
    wire _502;
    wire _503;
    wire _507;
    wire [64:0] _495;
    wire _496;
    wire _497;
    wire [64:0] _491;
    wire _493;
    wire _494;
    wire _498;
    wire _487;
    wire _488;
    wire [64:0] _483;
    wire [64:0] _482;
    wire _484;
    wire _485;
    wire _489;
    wire [64:0] _477;
    wire _478;
    wire _479;
    wire [64:0] _474;
    wire [64:0] _473;
    wire _475;
    wire _476;
    wire _480;
    wire [64:0] _468;
    wire _469;
    wire _470;
    wire [64:0] _465;
    wire [64:0] _464;
    wire _466;
    wire _467;
    wire _471;
    wire [64:0] _459;
    wire _460;
    wire _461;
    wire [64:0] _456;
    wire [64:0] _455;
    wire _457;
    wire _458;
    wire _462;
    wire [64:0] _450;
    wire _451;
    wire _452;
    wire [64:0] _447;
    wire [64:0] _446;
    wire _448;
    wire _449;
    wire _453;
    wire _442;
    wire _443;
    wire [64:0] _437;
    wire _439;
    wire _440;
    wire _444;
    wire [64:0] _432;
    wire _433;
    wire _434;
    wire [64:0] _429;
    wire [64:0] _428;
    wire _430;
    wire _431;
    wire _435;
    wire _424;
    wire _425;
    wire [64:0] _420;
    wire [64:0] _419;
    wire _421;
    wire _422;
    wire _426;
    wire _415;
    wire _416;
    wire [64:0] _410;
    wire _412;
    wire _413;
    wire _417;
    wire [64:0] _405;
    wire _406;
    wire _407;
    wire [64:0] _402;
    wire [64:0] _401;
    wire _403;
    wire _404;
    wire _408;
    wire [64:0] _396;
    wire _397;
    wire _398;
    wire [64:0] _392;
    wire _394;
    wire _395;
    wire _399;
    wire [64:0] _387;
    wire _388;
    wire _389;
    wire [64:0] _384;
    wire [64:0] _383;
    wire _385;
    wire _386;
    wire _390;
    wire [64:0] _378;
    wire _379;
    wire _380;
    wire [64:0] _374;
    wire _376;
    wire _377;
    wire _381;
    wire [64:0] _369;
    wire _370;
    wire _371;
    wire [64:0] _366;
    wire [64:0] _365;
    wire _367;
    wire _368;
    wire _372;
    wire [64:0] _360;
    wire _361;
    wire _362;
    wire [64:0] _357;
    wire [64:0] _356;
    wire _358;
    wire _359;
    wire _363;
    wire [64:0] _351;
    wire _352;
    wire _353;
    wire [64:0] _348;
    wire [64:0] _347;
    wire _349;
    wire _350;
    wire _354;
    wire [64:0] _342;
    wire _343;
    wire _344;
    wire [64:0] _339;
    wire [64:0] _338;
    wire _340;
    wire _341;
    wire _345;
    wire [64:0] _333;
    wire _334;
    wire _335;
    wire [64:0] _330;
    wire [64:0] _329;
    wire _331;
    wire _332;
    wire _336;
    wire _325;
    wire _326;
    wire [64:0] _320;
    wire _322;
    wire _323;
    wire _327;
    wire [64:0] _315;
    wire _316;
    wire _317;
    wire [64:0] _312;
    wire [64:0] _311;
    wire _313;
    wire _314;
    wire _318;
    wire _307;
    wire _308;
    wire [64:0] _303;
    wire [64:0] _302;
    wire _304;
    wire _305;
    wire _309;
    wire [64:0] _297;
    wire _298;
    wire _299;
    wire [64:0] _294;
    wire [64:0] _293;
    wire _295;
    wire _296;
    wire _300;
    wire [64:0] _288;
    wire _289;
    wire _290;
    wire [64:0] _285;
    wire [64:0] _284;
    wire _286;
    wire _287;
    wire _291;
    wire [64:0] _279;
    wire _280;
    wire _281;
    wire [64:0] _276;
    wire [64:0] _275;
    wire _277;
    wire _278;
    wire _282;
    wire [64:0] _270;
    wire _271;
    wire _272;
    wire [64:0] _267;
    wire [64:0] _266;
    wire _268;
    wire _269;
    wire _273;
    wire _262;
    wire _263;
    wire [64:0] _258;
    wire [64:0] _257;
    wire _259;
    wire _260;
    wire _264;
    wire _253;
    wire _254;
    wire [64:0] _249;
    wire [64:0] _248;
    wire _250;
    wire _251;
    wire _255;
    wire [64:0] _243;
    wire _244;
    wire _245;
    wire [64:0] _239;
    wire _241;
    wire _242;
    wire _246;
    wire [64:0] _234;
    wire _235;
    wire _236;
    wire [64:0] _231;
    wire [64:0] _230;
    wire _232;
    wire _233;
    wire _237;
    wire _226;
    wire _227;
    wire [64:0] _222;
    wire [64:0] _221;
    wire _223;
    wire _224;
    wire _228;
    wire [64:0] _216;
    wire _217;
    wire _218;
    wire [64:0] _213;
    wire [64:0] _212;
    wire _214;
    wire _215;
    wire _219;
    wire _208;
    wire _209;
    wire [64:0] _203;
    wire _205;
    wire _206;
    wire _210;
    wire [64:0] _198;
    wire _199;
    wire _200;
    wire [64:0] _194;
    wire _196;
    wire _197;
    wire _201;
    wire [64:0] _189;
    wire _190;
    wire _191;
    wire [64:0] _186;
    wire [64:0] _185;
    wire _187;
    wire _188;
    wire _192;
    wire [64:0] _180;
    wire _181;
    wire _182;
    wire [64:0] _177;
    wire [64:0] _176;
    wire _178;
    wire _179;
    wire _183;
    wire _172;
    wire _173;
    wire [64:0] _167;
    wire _169;
    wire _170;
    wire _174;
    wire [64:0] _162;
    wire _163;
    wire _164;
    wire [64:0] _159;
    wire [64:0] _158;
    wire _160;
    wire _161;
    wire _165;
    wire [64:0] _153;
    wire _154;
    wire _155;
    wire [64:0] _150;
    wire [64:0] _149;
    wire _151;
    wire _152;
    wire _156;
    wire _145;
    wire _146;
    wire [64:0] _140;
    wire _142;
    wire _143;
    wire _147;
    wire [64:0] _135;
    wire _136;
    wire _137;
    wire [64:0] _132;
    wire [64:0] _131;
    wire _133;
    wire _134;
    wire _138;
    wire [64:0] _126;
    wire _127;
    wire _128;
    wire [64:0] _122;
    wire _124;
    wire _125;
    wire _129;
    wire _118;
    wire _119;
    wire [64:0] _113;
    wire _115;
    wire _116;
    wire _120;
    wire [64:0] _108;
    wire _109;
    wire _110;
    wire [64:0] _105;
    wire [64:0] _104;
    wire _106;
    wire _107;
    wire _111;
    wire [64:0] _99;
    wire _100;
    wire _101;
    wire [64:0] _96;
    wire [64:0] _95;
    wire _97;
    wire _98;
    wire _102;
    wire _91;
    wire _92;
    wire [64:0] _86;
    wire _88;
    wire _89;
    wire _93;
    wire [64:0] _81;
    wire _82;
    wire _83;
    wire [64:0] _78;
    wire [64:0] _77;
    wire _79;
    wire _80;
    wire _84;
    wire [64:0] _72;
    wire _73;
    wire _74;
    wire [64:0] _69;
    wire [64:0] _68;
    wire _70;
    wire _71;
    wire _75;
    wire [64:0] _63;
    wire _64;
    wire _65;
    wire [64:0] _59;
    wire _61;
    wire _62;
    wire _66;
    wire _55;
    wire _56;
    wire [64:0] _50;
    wire _52;
    wire _53;
    wire _57;
    wire _46;
    wire _47;
    wire [64:0] _42;
    wire [64:0] _41;
    wire _43;
    wire _44;
    wire _48;
    wire [64:0] _36;
    wire _37;
    wire _38;
    wire [64:0] _33;
    wire [64:0] _32;
    wire _34;
    wire _35;
    wire _39;
    wire _28;
    wire _29;
    wire [64:0] _24;
    wire [64:0] _23;
    wire _25;
    wire _26;
    wire _30;
    wire [64:0] _19;
    wire _20;
    wire _21;
    wire [64:0] _16;
    wire [63:0] _10;
    wire gnd;
    wire [64:0] _15;
    wire _17;
    wire _18;
    wire _22;
    wire _31;
    wire _40;
    wire _49;
    wire _58;
    wire _67;
    wire _76;
    wire _85;
    wire _94;
    wire _103;
    wire _112;
    wire _121;
    wire _130;
    wire _139;
    wire _148;
    wire _157;
    wire _166;
    wire _175;
    wire _184;
    wire _193;
    wire _202;
    wire _211;
    wire _220;
    wire _229;
    wire _238;
    wire _247;
    wire _256;
    wire _265;
    wire _274;
    wire _283;
    wire _292;
    wire _301;
    wire _310;
    wire _319;
    wire _328;
    wire _337;
    wire _346;
    wire _355;
    wire _364;
    wire _373;
    wire _382;
    wire _391;
    wire _400;
    wire _409;
    wire _418;
    wire _427;
    wire _436;
    wire _445;
    wire _454;
    wire _463;
    wire _472;
    wire _481;
    wire _490;
    wire _499;
    wire _508;
    wire _517;
    wire _526;
    wire _535;
    wire _544;
    wire _553;
    wire _562;
    wire _571;
    wire _580;
    wire _589;
    wire _598;
    wire _607;
    wire _616;
    wire _625;
    wire _634;
    wire _643;
    wire _652;
    wire _661;
    wire _670;
    wire _679;
    wire _688;
    wire _697;
    wire _706;
    wire _715;
    wire _724;
    wire _733;
    wire _742;
    wire _751;
    wire _760;
    wire _769;
    wire _778;
    wire _787;
    wire _796;
    wire _805;
    wire _814;
    wire _823;
    wire _832;
    wire _841;
    wire _850;
    wire _859;
    wire _868;
    wire _877;
    wire _886;
    wire _895;
    wire _904;
    wire _913;
    wire _922;
    wire _931;
    wire _940;
    wire _949;
    wire _958;
    wire _967;
    wire _976;
    wire _985;
    wire _994;
    wire _1003;
    wire _1012;
    wire _1021;
    wire _1030;
    wire _1039;
    wire _1048;
    wire _1057;
    wire _1066;
    wire _1075;
    wire _1084;
    wire _1093;
    wire _1102;
    wire _1111;
    wire _1120;
    wire _1129;
    wire _1138;
    wire _1147;
    wire _1156;
    wire _1165;
    wire _1174;
    wire _1183;
    wire _1192;
    wire _1201;
    wire _1210;
    wire _1219;
    wire _1228;
    wire _1237;
    wire _1246;
    wire _1255;
    wire _1264;
    wire _1273;
    wire _1282;
    wire _1291;
    wire _1300;
    wire _1309;
    wire _1318;
    wire _1327;
    wire _1336;
    wire _1345;
    wire _1354;
    wire _1363;
    wire _1372;
    wire _1381;
    wire _1390;
    wire _1399;
    wire _1408;
    wire _1417;
    wire _1426;
    wire _1435;
    wire _1444;
    wire _1453;
    wire _1462;
    wire _1471;
    wire _1480;
    wire _1489;
    wire _1498;
    wire _1507;
    wire _1516;
    wire _1525;
    wire _1534;
    wire _1543;
    wire _1552;
    wire _1561;
    wire _1570;
    wire _1579;
    wire _1588;
    wire _1597;
    wire _1606;
    wire _1615;
    wire _1624;
    wire _1633;
    wire _1642;
    wire _1651;
    wire _1660;
    wire _1669;
    wire _1678;
    wire _1687;
    wire _1696;
    assign _2 = valid;
    assign _1697 = _1696 & _2;
    assign _13 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _4 = clear;
    assign _6 = clock;
    assign _1699 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    assign _1700 = _1698 + _1699;
    assign _7 = _1700;
    always @(posedge _6) begin
        if (_4)
            _1698 <= _13;
        else
            if (_1697)
                _1698 <= _7;
    end
    assign _1692 = 65'b00000000000000000110101011010010001001110000000001000101101000000;
    assign _1693 = _1692 < _1688;
    assign _1694 = ~ _1693;
    assign _1689 = 65'b00000000000000000110100111010010010011100010111011000001111111011;
    assign _1688 = { gnd,
                     _10 };
    assign _1690 = _1688 < _1689;
    assign _1691 = ~ _1690;
    assign _1695 = _1691 & _1694;
    assign _1683 = 65'b00000000000000001000011110101000111001101010101110001100000110111;
    assign _1684 = _1683 < _1679;
    assign _1685 = ~ _1684;
    assign _1680 = 65'b00000000000000001000010100001101111001111111000010111010010111110;
    assign _1679 = { gnd,
                     _10 };
    assign _1681 = _1679 < _1680;
    assign _1682 = ~ _1681;
    assign _1686 = _1682 & _1685;
    assign _1674 = 65'b00000000000000000100010110110100111101111010010010100111101111000;
    assign _1675 = _1674 < _1670;
    assign _1676 = ~ _1675;
    assign _1671 = 65'b00000000000000000100010100011111001111111100010011111001011101001;
    assign _1670 = { gnd,
                     _10 };
    assign _1672 = _1670 < _1671;
    assign _1673 = ~ _1672;
    assign _1677 = _1673 & _1676;
    assign _1665 = 65'b00000000000000000001000001100110010010011101001111110110111010101;
    assign _1666 = _1665 < _1661;
    assign _1667 = ~ _1666;
    assign _1662 = 65'b00000000000000000000111110101001011010010010100101000001110001000;
    assign _1661 = { gnd,
                     _10 };
    assign _1663 = _1661 < _1662;
    assign _1664 = ~ _1663;
    assign _1668 = _1664 & _1667;
    assign _1656 = 65'b00000000000000001010100010110011010111001100000010010100100010100;
    assign _1657 = _1656 < _1652;
    assign _1658 = ~ _1657;
    assign _1653 = 65'b00000000000000001010011001010000111110010110111101101100000000110;
    assign _1652 = { gnd,
                     _10 };
    assign _1654 = _1652 < _1653;
    assign _1655 = ~ _1654;
    assign _1659 = _1655 & _1658;
    assign _1647 = 65'b00000000000000000010111001110101010000001101101110111111100101100;
    assign _1648 = _1647 < _1643;
    assign _1649 = ~ _1648;
    assign _1644 = 65'b00000000000000000010111001001110110011001010001111001000000010010;
    assign _1643 = { gnd,
                     _10 };
    assign _1645 = _1643 < _1644;
    assign _1646 = ~ _1645;
    assign _1650 = _1646 & _1649;
    assign _1638 = 65'b00000000000000001100110010001010100011000111001101110100100100001;
    assign _1639 = _1638 < _1634;
    assign _1640 = ~ _1639;
    assign _1635 = 65'b00000000000000001100101001000110101010010010110101001100111110100;
    assign _1634 = { gnd,
                     _10 };
    assign _1636 = _1634 < _1635;
    assign _1637 = ~ _1636;
    assign _1641 = _1637 & _1640;
    assign _1629 = 65'b00000000000000000011101001110110011000111011000110101110001100100;
    assign _1630 = _1629 < _1625;
    assign _1631 = ~ _1630;
    assign _1626 = 65'b00000000000000000011100000011000010001011011010011001001010111110;
    assign _1625 = { gnd,
                     _10 };
    assign _1627 = _1625 < _1626;
    assign _1628 = ~ _1627;
    assign _1632 = _1628 & _1631;
    assign _1620 = 65'b00000000000000001111111001001000010100011010100000010110000001101;
    assign _1621 = _1620 < _1616;
    assign _1622 = ~ _1621;
    assign _1617 = 65'b00000000000000001111110001010000000010000111100001000010011010111;
    assign _1616 = { gnd,
                     _10 };
    assign _1618 = _1616 < _1617;
    assign _1619 = ~ _1618;
    assign _1623 = _1619 & _1622;
    assign _1611 = 65'b00000000000000000111101010101001011010010000011101001000100001011;
    assign _1612 = _1611 < _1607;
    assign _1613 = ~ _1612;
    assign _1608 = 65'b00000000000000000111011100101001011100011011011110111001101001011;
    assign _1607 = { gnd,
                     _10 };
    assign _1609 = _1607 < _1608;
    assign _1610 = ~ _1609;
    assign _1614 = _1610 & _1613;
    assign _1602 = 65'b00000000000000000100111101111110000001111101101000000100111111111;
    assign _1603 = _1602 < _1598;
    assign _1604 = ~ _1603;
    assign _1599 = 65'b00000000000000000100111100100101001000010111101101000110110111111;
    assign _1598 = { gnd,
                     _10 };
    assign _1600 = _1598 < _1599;
    assign _1601 = ~ _1600;
    assign _1605 = _1601 & _1604;
    assign _1593 = 65'b00000000000000000101000111000001110111101000110000110111100100110;
    assign _1594 = _1593 < _1589;
    assign _1595 = ~ _1594;
    assign _1590 = 65'b00000000000000000101000110001010000011101010100010000111111100000;
    assign _1589 = { gnd,
                     _10 };
    assign _1591 = _1589 < _1590;
    assign _1592 = ~ _1591;
    assign _1596 = _1592 & _1595;
    assign _1584 = 65'b00000000000000000100100100011101100000011111100101001101001000001;
    assign _1585 = _1584 < _1580;
    assign _1586 = ~ _1585;
    assign _1581 = 65'b00000000000000000100100001111100000100101111110111111001000011001;
    assign _1580 = { gnd,
                     _10 };
    assign _1582 = _1580 < _1581;
    assign _1583 = ~ _1582;
    assign _1587 = _1583 & _1586;
    assign _1575 = 65'b00000000000000000110100001100010001111110010001000100010010100010;
    assign _1576 = _1575 < _1571;
    assign _1577 = ~ _1576;
    assign _1572 = 65'b00000000000000000110010011100000010110101110100011100000001001010;
    assign _1571 = { gnd,
                     _10 };
    assign _1573 = _1571 < _1572;
    assign _1574 = ~ _1573;
    assign _1578 = _1574 & _1577;
    assign _1566 = 65'b00000000000000000101101011001110101000100001010111011000110110101;
    assign _1567 = _1566 < _1562;
    assign _1568 = ~ _1567;
    assign _1562 = { gnd,
                     _10 };
    assign _1564 = _1562 < _1566;
    assign _1565 = ~ _1564;
    assign _1569 = _1565 & _1568;
    assign _1557 = 65'b00000000000000001101100011000010010001011110011101001001110110101;
    assign _1558 = _1557 < _1553;
    assign _1559 = ~ _1558;
    assign _1554 = 65'b00000000000000001101100000100010100000100000010010010111111000011;
    assign _1553 = { gnd,
                     _10 };
    assign _1555 = _1553 < _1554;
    assign _1556 = ~ _1555;
    assign _1560 = _1556 & _1559;
    assign _1548 = 65'b00000000000000000100010100111101011010000100111010010011000110110;
    assign _1549 = _1548 < _1544;
    assign _1550 = ~ _1549;
    assign _1545 = 65'b00000000000000000100010010111001111011110010010110011000001011100;
    assign _1544 = { gnd,
                     _10 };
    assign _1546 = _1544 < _1545;
    assign _1547 = ~ _1546;
    assign _1551 = _1547 & _1550;
    assign _1539 = 65'b00000000000000000101011010000111111110000100011011110010000100110;
    assign _1540 = _1539 < _1535;
    assign _1541 = ~ _1540;
    assign _1536 = 65'b00000000000000000101001100100011001101110100100010000000011000011;
    assign _1535 = { gnd,
                     _10 };
    assign _1537 = _1535 < _1536;
    assign _1538 = ~ _1537;
    assign _1542 = _1538 & _1541;
    assign _1530 = 65'b00000000000000000100111010101111101101100101100010011110011001000;
    assign _1531 = _1530 < _1526;
    assign _1532 = ~ _1531;
    assign _1527 = 65'b00000000000000000100111001010001011100011011001111011111111110011;
    assign _1526 = { gnd,
                     _10 };
    assign _1528 = _1526 < _1527;
    assign _1529 = ~ _1528;
    assign _1533 = _1529 & _1532;
    assign _1521 = 65'b00000000000000000110110011010111000100011100101000110001000101111;
    assign _1522 = _1521 < _1517;
    assign _1523 = ~ _1522;
    assign _1517 = { gnd,
                     _10 };
    assign _1519 = _1517 < _1689;
    assign _1520 = ~ _1519;
    assign _1524 = _1520 & _1523;
    assign _1512 = 65'b00000000000000000101110101010111100010101101011010010111010000101;
    assign _1513 = _1512 < _1508;
    assign _1514 = ~ _1513;
    assign _1509 = 65'b00000000000000000101110001011100101100111000100101010010111010101;
    assign _1508 = { gnd,
                     _10 };
    assign _1510 = _1508 < _1509;
    assign _1511 = ~ _1510;
    assign _1515 = _1511 & _1514;
    assign _1503 = 65'b00000000000000001011010110111110010101001010011010011100001000100;
    assign _1504 = _1503 < _1499;
    assign _1505 = ~ _1504;
    assign _1500 = 65'b00000000000000001011001010001010111011110001100010101001100001011;
    assign _1499 = { gnd,
                     _10 };
    assign _1501 = _1499 < _1500;
    assign _1502 = ~ _1501;
    assign _1506 = _1502 & _1505;
    assign _1494 = 65'b00000000000000000010110011110110010101100000101101010000010001001;
    assign _1495 = _1494 < _1490;
    assign _1496 = ~ _1495;
    assign _1491 = 65'b00000000000000000010101011111100100000110011100001011110011011101;
    assign _1490 = { gnd,
                     _10 };
    assign _1492 = _1490 < _1491;
    assign _1493 = ~ _1492;
    assign _1497 = _1493 & _1496;
    assign _1485 = 65'b00000000000000001001011001011001101010001101110001111011011111001;
    assign _1486 = _1485 < _1481;
    assign _1487 = ~ _1486;
    assign _1482 = 65'b00000000000000001001011000111100100001110001011000000101011101000;
    assign _1481 = { gnd,
                     _10 };
    assign _1483 = _1481 < _1482;
    assign _1484 = ~ _1483;
    assign _1488 = _1484 & _1487;
    assign _1476 = 65'b00000000000000001101111000000111101100111001000011111111110111111;
    assign _1477 = _1476 < _1472;
    assign _1478 = ~ _1477;
    assign _1473 = 65'b00000000000000001101110111010000010110001001101101001100101101111;
    assign _1472 = { gnd,
                     _10 };
    assign _1474 = _1472 < _1473;
    assign _1475 = ~ _1474;
    assign _1479 = _1475 & _1478;
    assign _1467 = 65'b00000000000000001001100001111011100010100011101100000100101000111;
    assign _1468 = _1467 < _1463;
    assign _1469 = ~ _1468;
    assign _1464 = 65'b00000000000000001001011111010010001101101000001111011011001100000;
    assign _1463 = { gnd,
                     _10 };
    assign _1465 = _1463 < _1464;
    assign _1466 = ~ _1465;
    assign _1470 = _1466 & _1469;
    assign _1458 = 65'b00000000000000001101100000010010110001011000011001000111001110100;
    assign _1459 = _1458 < _1454;
    assign _1460 = ~ _1459;
    assign _1455 = 65'b00000000000000001101011101001101111101010110110111010100101001011;
    assign _1454 = { gnd,
                     _10 };
    assign _1456 = _1454 < _1455;
    assign _1457 = ~ _1456;
    assign _1461 = _1457 & _1460;
    assign _1449 = 65'b00000000000000000100011101011100110010001010011101010001000111010;
    assign _1450 = _1449 < _1445;
    assign _1451 = ~ _1450;
    assign _1446 = 65'b00000000000000000100011011010000011100010100100110111101011010110;
    assign _1445 = { gnd,
                     _10 };
    assign _1447 = _1445 < _1446;
    assign _1448 = ~ _1447;
    assign _1452 = _1448 & _1451;
    assign _1440 = 65'b00000000000000000100111011100010000110010101011010000010000101111;
    assign _1441 = _1440 < _1436;
    assign _1442 = ~ _1441;
    assign _1437 = 65'b00000000000000000100111011001010110010010010001111010001010000100;
    assign _1436 = { gnd,
                     _10 };
    assign _1438 = _1436 < _1437;
    assign _1439 = ~ _1438;
    assign _1443 = _1439 & _1442;
    assign _1431 = 65'b00000000000000001101010010011001010011110000010010001110000111001;
    assign _1432 = _1431 < _1427;
    assign _1433 = ~ _1432;
    assign _1428 = 65'b00000000000000001101001100010100010110100010000111111110010100100;
    assign _1427 = { gnd,
                     _10 };
    assign _1429 = _1427 < _1428;
    assign _1430 = ~ _1429;
    assign _1434 = _1430 & _1433;
    assign _1423 = _1473 < _1418;
    assign _1424 = ~ _1423;
    assign _1419 = 65'b00000000000000001101110101110010010101011000110100100110101100011;
    assign _1418 = { gnd,
                     _10 };
    assign _1420 = _1418 < _1419;
    assign _1421 = ~ _1420;
    assign _1425 = _1421 & _1424;
    assign _1413 = 65'b00000000000000001011101010000011111010100011000011100111100110000;
    assign _1414 = _1413 < _1409;
    assign _1415 = ~ _1414;
    assign _1409 = { gnd,
                     _10 };
    assign _1411 = _1409 < _1413;
    assign _1412 = ~ _1411;
    assign _1416 = _1412 & _1415;
    assign _1404 = 65'b00000000000000001111100101100110010011101101111001111001011100010;
    assign _1405 = _1404 < _1400;
    assign _1406 = ~ _1405;
    assign _1401 = 65'b00000000000000001111100011100101111001101111010011001010101001101;
    assign _1400 = { gnd,
                     _10 };
    assign _1402 = _1400 < _1401;
    assign _1403 = ~ _1402;
    assign _1407 = _1403 & _1406;
    assign _1395 = 65'b00000000000000001010101111110100000011000100111011011001100011101;
    assign _1396 = _1395 < _1391;
    assign _1397 = ~ _1396;
    assign _1391 = { gnd,
                     _10 };
    assign _1393 = _1391 < _1395;
    assign _1394 = ~ _1393;
    assign _1398 = _1394 & _1397;
    assign _1386 = 65'b00000000000000000011000010000010011111110011100010101001101110110;
    assign _1387 = _1386 < _1382;
    assign _1388 = ~ _1387;
    assign _1383 = 65'b00000000000000000011000001001010000110001111100000100111110111111;
    assign _1382 = { gnd,
                     _10 };
    assign _1384 = _1382 < _1383;
    assign _1385 = ~ _1384;
    assign _1389 = _1385 & _1388;
    assign _1377 = 65'b00000000000000000010011111001011101111110101000001111010001001011;
    assign _1378 = _1377 < _1373;
    assign _1379 = ~ _1378;
    assign _1374 = 65'b00000000000000000010011001101100110001101001110110000100100101010;
    assign _1373 = { gnd,
                     _10 };
    assign _1375 = _1373 < _1374;
    assign _1376 = ~ _1375;
    assign _1380 = _1376 & _1379;
    assign _1368 = 65'b00000000000000000001001000111011001111001011110111110110011101101;
    assign _1369 = _1368 < _1364;
    assign _1370 = ~ _1369;
    assign _1365 = 65'b00000000000000000001000101101100100101110001010010110100000001110;
    assign _1364 = { gnd,
                     _10 };
    assign _1366 = _1364 < _1365;
    assign _1367 = ~ _1366;
    assign _1371 = _1367 & _1370;
    assign _1359 = 65'b00000000000000000100111000101000001110000000110110010111101100100;
    assign _1360 = _1359 < _1355;
    assign _1361 = ~ _1360;
    assign _1356 = 65'b00000000000000000100110111100010010101110100111010110110101100010;
    assign _1355 = { gnd,
                     _10 };
    assign _1357 = _1355 < _1356;
    assign _1358 = ~ _1357;
    assign _1362 = _1358 & _1361;
    assign _1350 = 65'b00000000000000001001100000001111111111011111101111001101110011110;
    assign _1351 = _1350 < _1346;
    assign _1352 = ~ _1351;
    assign _1347 = 65'b00000000000000001001011101010111011010011110011110100100111111001;
    assign _1346 = { gnd,
                     _10 };
    assign _1348 = _1346 < _1347;
    assign _1349 = ~ _1348;
    assign _1353 = _1349 & _1352;
    assign _1341 = 65'b00000000000000000001101000001010011010011000001101111101111101110;
    assign _1342 = _1341 < _1337;
    assign _1343 = ~ _1342;
    assign _1337 = { gnd,
                     _10 };
    assign _1339 = _1337 < _1341;
    assign _1340 = ~ _1339;
    assign _1344 = _1340 & _1343;
    assign _1332 = 65'b00000000000000000010001010100001011011001010101000100000000101111;
    assign _1333 = _1332 < _1328;
    assign _1334 = ~ _1333;
    assign _1329 = 65'b00000000000000000010000000101011111111110011101100001100011011111;
    assign _1328 = { gnd,
                     _10 };
    assign _1330 = _1328 < _1329;
    assign _1331 = ~ _1330;
    assign _1335 = _1331 & _1334;
    assign _1323 = 65'b00000000000000000010111100000101001111110001111010011101111100111;
    assign _1324 = _1323 < _1319;
    assign _1325 = ~ _1324;
    assign _1320 = 65'b00000000000000000010111011101100000110111110111100000100001000010;
    assign _1319 = { gnd,
                     _10 };
    assign _1321 = _1319 < _1320;
    assign _1322 = ~ _1321;
    assign _1326 = _1322 & _1325;
    assign _1314 = 65'b00000000000000000100011010000111000101100100111111001101011000100;
    assign _1315 = _1314 < _1310;
    assign _1316 = ~ _1315;
    assign _1311 = 65'b00000000000000000100010111010110110101001110101011101010010001011;
    assign _1310 = { gnd,
                     _10 };
    assign _1312 = _1310 < _1311;
    assign _1313 = ~ _1312;
    assign _1317 = _1313 & _1316;
    assign _1305 = 65'b00000000000000001001100110110000110110001100100100111011101000101;
    assign _1306 = _1305 < _1301;
    assign _1307 = ~ _1306;
    assign _1302 = 65'b00000000000000001001100100000110101001010111000100111000011000011;
    assign _1301 = { gnd,
                     _10 };
    assign _1303 = _1301 < _1302;
    assign _1304 = ~ _1303;
    assign _1308 = _1304 & _1307;
    assign _1297 = _1566 < _1292;
    assign _1298 = ~ _1297;
    assign _1293 = 65'b00000000000000000101011100101110110110000100000100111000100010000;
    assign _1292 = { gnd,
                     _10 };
    assign _1294 = _1292 < _1293;
    assign _1295 = ~ _1294;
    assign _1299 = _1295 & _1298;
    assign _1287 = 65'b00000000000000000100111101001000100011001010000100111110100001010;
    assign _1288 = _1287 < _1283;
    assign _1289 = ~ _1288;
    assign _1283 = { gnd,
                     _10 };
    assign _1285 = _1283 < _1599;
    assign _1286 = ~ _1285;
    assign _1290 = _1286 & _1289;
    assign _1278 = 65'b00000000000000001001000111000001101011101001000101100110011101011;
    assign _1279 = _1278 < _1274;
    assign _1280 = ~ _1279;
    assign _1275 = 65'b00000000000000001000111010111100110111011110001110011100011111111;
    assign _1274 = { gnd,
                     _10 };
    assign _1276 = _1274 < _1275;
    assign _1277 = ~ _1276;
    assign _1281 = _1277 & _1280;
    assign _1269 = 65'b00000000000000000111011001000100110001110101000110001110010001010;
    assign _1270 = _1269 < _1265;
    assign _1271 = ~ _1270;
    assign _1265 = { gnd,
                     _10 };
    assign _1267 = _1265 < _1269;
    assign _1268 = ~ _1267;
    assign _1272 = _1268 & _1271;
    assign _1260 = 65'b00000000000000001100001010110111011001011010101000101101100010101;
    assign _1261 = _1260 < _1256;
    assign _1262 = ~ _1261;
    assign _1256 = { gnd,
                     _10 };
    assign _1258 = _1256 < _1260;
    assign _1259 = ~ _1258;
    assign _1263 = _1259 & _1262;
    assign _1251 = 65'b00000000000000001101111110110000111111111011001100001100010110001;
    assign _1252 = _1251 < _1247;
    assign _1253 = ~ _1252;
    assign _1248 = 65'b00000000000000001101111110000101110001000111000011000110001000100;
    assign _1247 = { gnd,
                     _10 };
    assign _1249 = _1247 < _1248;
    assign _1250 = ~ _1249;
    assign _1254 = _1250 & _1253;
    assign _1242 = 65'b00000000000000000011000000110110110111101001110000001110011010010;
    assign _1243 = _1242 < _1238;
    assign _1244 = ~ _1243;
    assign _1239 = 65'b00000000000000000010111111101111001100000011101100100010111000110;
    assign _1238 = { gnd,
                     _10 };
    assign _1240 = _1238 < _1239;
    assign _1241 = ~ _1240;
    assign _1245 = _1241 & _1244;
    assign _1233 = 65'b00000000000000000010011001101100110001101001110110000100100101000;
    assign _1234 = _1233 < _1229;
    assign _1235 = ~ _1234;
    assign _1230 = 65'b00000000000000000010010100010100111001101110111001111110001100000;
    assign _1229 = { gnd,
                     _10 };
    assign _1231 = _1229 < _1230;
    assign _1232 = ~ _1231;
    assign _1236 = _1232 & _1235;
    assign _1224 = 65'b00000000000000001011000101111101000001100101111100111001010101000;
    assign _1225 = _1224 < _1220;
    assign _1226 = ~ _1225;
    assign _1221 = 65'b00000000000000001010111000100101011110111101011111110000111100101;
    assign _1220 = { gnd,
                     _10 };
    assign _1222 = _1220 < _1221;
    assign _1223 = ~ _1222;
    assign _1227 = _1223 & _1226;
    assign _1215 = 65'b00000000000000000011010110111100110001111101111110100010111100111;
    assign _1216 = _1215 < _1211;
    assign _1217 = ~ _1216;
    assign _1212 = 65'b00000000000000000011001101111000011001111101001000110100100110001;
    assign _1211 = { gnd,
                     _10 };
    assign _1213 = _1211 < _1212;
    assign _1214 = ~ _1213;
    assign _1218 = _1214 & _1217;
    assign _1206 = 65'b00000000000000001111111110011100110011010100100110001010010101111;
    assign _1207 = _1206 < _1202;
    assign _1208 = ~ _1207;
    assign _1203 = 65'b00000000000000001111111001001000010100011010100000010110000001111;
    assign _1202 = { gnd,
                     _10 };
    assign _1204 = _1202 < _1203;
    assign _1205 = ~ _1204;
    assign _1209 = _1205 & _1208;
    assign _1198 = _1287 < _1193;
    assign _1199 = ~ _1198;
    assign _1193 = { gnd,
                     _10 };
    assign _1195 = _1193 < _1599;
    assign _1196 = ~ _1195;
    assign _1200 = _1196 & _1199;
    assign _1188 = 65'b00000000000000001101101000011110000010001101001110010010000001000;
    assign _1189 = _1188 < _1184;
    assign _1190 = ~ _1189;
    assign _1185 = 65'b00000000000000001101100101110111111010010101010010110101000010011;
    assign _1184 = { gnd,
                     _10 };
    assign _1186 = _1184 < _1185;
    assign _1187 = ~ _1186;
    assign _1191 = _1187 & _1190;
    assign _1179 = 65'b00000000000000001110100001010111110111110100010110101100000100110;
    assign _1180 = _1179 < _1175;
    assign _1181 = ~ _1180;
    assign _1175 = { gnd,
                     _10 };
    assign _1177 = _1175 < _1179;
    assign _1178 = ~ _1177;
    assign _1182 = _1178 & _1181;
    assign _1170 = 65'b00000000000000001010101111110100000011000100111011011001100011100;
    assign _1171 = _1170 < _1166;
    assign _1172 = ~ _1171;
    assign _1167 = 65'b00000000000000001010101010000101010011011111111010100100010100101;
    assign _1166 = { gnd,
                     _10 };
    assign _1168 = _1166 < _1167;
    assign _1169 = ~ _1168;
    assign _1173 = _1169 & _1172;
    assign _1161 = 65'b00000000000000000000110000001111000011000001001010101100110110011;
    assign _1162 = _1161 < _1157;
    assign _1163 = ~ _1162;
    assign _1158 = 65'b00000000000000000000101100101010010000101100001100001011001010000;
    assign _1157 = { gnd,
                     _10 };
    assign _1159 = _1157 < _1158;
    assign _1160 = ~ _1159;
    assign _1164 = _1160 & _1163;
    assign _1152 = 65'b00000000000000001101000111100010001111010101000100100001000111100;
    assign _1153 = _1152 < _1148;
    assign _1154 = ~ _1153;
    assign _1149 = 65'b00000000000000001100111000100111110011010100111111010111110110110;
    assign _1148 = { gnd,
                     _10 };
    assign _1150 = _1148 < _1149;
    assign _1151 = ~ _1150;
    assign _1155 = _1151 & _1154;
    assign _1143 = 65'b00000000000000001001101011100110001001011000101011111111011101110;
    assign _1144 = _1143 < _1139;
    assign _1145 = ~ _1144;
    assign _1140 = 65'b00000000000000001001101001001000101000100101111000100111110001011;
    assign _1139 = { gnd,
                     _10 };
    assign _1141 = _1139 < _1140;
    assign _1142 = ~ _1141;
    assign _1146 = _1142 & _1145;
    assign _1134 = 65'b00000000000000000000100000110101000111101100011111000111010000100;
    assign _1135 = _1134 < _1130;
    assign _1136 = ~ _1135;
    assign _1131 = 65'b00000000000000000000010011110111100010101000101011110011100011010;
    assign _1130 = { gnd,
                     _10 };
    assign _1132 = _1130 < _1131;
    assign _1133 = ~ _1132;
    assign _1137 = _1133 & _1136;
    assign _1125 = 65'b00000000000000001001010100010101011111000010110100101000110010110;
    assign _1126 = _1125 < _1121;
    assign _1127 = ~ _1126;
    assign _1122 = 65'b00000000000000001001010011010000100110010011011000011000101010101;
    assign _1121 = { gnd,
                     _10 };
    assign _1123 = _1121 < _1122;
    assign _1124 = ~ _1123;
    assign _1128 = _1124 & _1127;
    assign _1116 = 65'b00000000000000000100001100000110100110110111000010000011000110001;
    assign _1117 = _1116 < _1112;
    assign _1118 = ~ _1117;
    assign _1113 = 65'b00000000000000000100000010001000011000101101110111000111101100010;
    assign _1112 = { gnd,
                     _10 };
    assign _1114 = _1112 < _1113;
    assign _1115 = ~ _1114;
    assign _1119 = _1115 & _1118;
    assign _1107 = 65'b00000000000000001001110111000111111110011011111111010000111101000;
    assign _1108 = _1107 < _1103;
    assign _1109 = ~ _1108;
    assign _1104 = 65'b00000000000000001001110000000001011001010101001000001000001010101;
    assign _1103 = { gnd,
                     _10 };
    assign _1105 = _1103 < _1104;
    assign _1106 = ~ _1105;
    assign _1110 = _1106 & _1109;
    assign _1098 = 65'b00000000000000001001011000011000010010010011101011110100001010000;
    assign _1099 = _1098 < _1094;
    assign _1100 = ~ _1099;
    assign _1095 = 65'b00000000000000001001010111111110110111100010010111000010000000101;
    assign _1094 = { gnd,
                     _10 };
    assign _1096 = _1094 < _1095;
    assign _1097 = ~ _1096;
    assign _1101 = _1097 & _1100;
    assign _1089 = 65'b00000000000000001101101111010110000010001000001111000100111101111;
    assign _1090 = _1089 < _1085;
    assign _1091 = ~ _1090;
    assign _1086 = 65'b00000000000000001101101101110001111011011110110000111100111010100;
    assign _1085 = { gnd,
                     _10 };
    assign _1087 = _1085 < _1086;
    assign _1088 = ~ _1087;
    assign _1092 = _1088 & _1091;
    assign _1080 = 65'b00000000000000000001000100101110000110101110000110101100101101011;
    assign _1081 = _1080 < _1076;
    assign _1082 = ~ _1081;
    assign _1077 = 65'b00000000000000000001000010010111100010001000001110001101111110110;
    assign _1076 = { gnd,
                     _10 };
    assign _1078 = _1076 < _1077;
    assign _1079 = ~ _1078;
    assign _1083 = _1079 & _1082;
    assign _1071 = 65'b00000000000000001001010110101101011011001010000101101001000000011;
    assign _1072 = _1071 < _1067;
    assign _1073 = ~ _1072;
    assign _1068 = 65'b00000000000000001001010101001011000101001110010100000111000011101;
    assign _1067 = { gnd,
                     _10 };
    assign _1069 = _1067 < _1068;
    assign _1070 = ~ _1069;
    assign _1074 = _1070 & _1073;
    assign _1062 = 65'b00000000000000001001001011001111010101001100110011001000000110110;
    assign _1063 = _1062 < _1058;
    assign _1064 = ~ _1063;
    assign _1059 = 65'b00000000000000001001001010001001000010001001101000001110011100001;
    assign _1058 = { gnd,
                     _10 };
    assign _1060 = _1058 < _1059;
    assign _1061 = ~ _1060;
    assign _1065 = _1061 & _1064;
    assign _1054 = _1359 < _1049;
    assign _1055 = ~ _1054;
    assign _1049 = { gnd,
                     _10 };
    assign _1051 = _1049 < _1356;
    assign _1052 = ~ _1051;
    assign _1056 = _1052 & _1055;
    assign _1044 = 65'b00000000000000001001100101001000100000101011110101111011011101000;
    assign _1045 = _1044 < _1040;
    assign _1046 = ~ _1045;
    assign _1041 = 65'b00000000000000001001100010011010010011001110001100000000110101011;
    assign _1040 = { gnd,
                     _10 };
    assign _1042 = _1040 < _1041;
    assign _1043 = ~ _1042;
    assign _1047 = _1043 & _1046;
    assign _1035 = 65'b00000000000000001001101101100101010011101011100111100010001001010;
    assign _1036 = _1035 < _1031;
    assign _1037 = ~ _1036;
    assign _1032 = 65'b00000000000000001001101010110110010111111001001001011100001100011;
    assign _1031 = { gnd,
                     _10 };
    assign _1033 = _1031 < _1032;
    assign _1034 = ~ _1033;
    assign _1038 = _1034 & _1037;
    assign _1026 = 65'b00000000000000001101101101010100000110011110100000010111111000001;
    assign _1027 = _1026 < _1022;
    assign _1028 = ~ _1027;
    assign _1023 = 65'b00000000000000001101101010110110110010010111110110111001010101010;
    assign _1022 = { gnd,
                     _10 };
    assign _1024 = _1022 < _1023;
    assign _1025 = ~ _1024;
    assign _1029 = _1025 & _1028;
    assign _1018 = _1638 < _1013;
    assign _1019 = ~ _1018;
    assign _1014 = 65'b00000000000000001100101100000111101000110101100001011011101111100;
    assign _1013 = { gnd,
                     _10 };
    assign _1015 = _1013 < _1014;
    assign _1016 = ~ _1015;
    assign _1020 = _1016 & _1019;
    assign _1008 = 65'b00000000000000000000111010000101101000000010110111000111001000100;
    assign _1009 = _1008 < _1004;
    assign _1010 = ~ _1009;
    assign _1005 = 65'b00000000000000000000110111100000101101100110111000000010101001011;
    assign _1004 = { gnd,
                     _10 };
    assign _1006 = _1004 < _1005;
    assign _1007 = ~ _1006;
    assign _1011 = _1007 & _1010;
    assign _999 = 65'b00000000000000000111111011010100000110001101001101011111011110101;
    assign _1000 = _999 < _995;
    assign _1001 = ~ _1000;
    assign _996 = 65'b00000000000000000111101111111110001101101101110010001101100011011;
    assign _995 = { gnd,
                    _10 };
    assign _997 = _995 < _996;
    assign _998 = ~ _997;
    assign _1002 = _998 & _1001;
    assign _990 = 65'b00000000000000001010111000100101011110111101011111110000111100100;
    assign _991 = _990 < _986;
    assign _992 = ~ _991;
    assign _986 = { gnd,
                    _10 };
    assign _988 = _986 < _990;
    assign _989 = ~ _988;
    assign _993 = _989 & _992;
    assign _981 = 65'b00000000000000001101110000001010100111110110011111101011011000000;
    assign _982 = _981 < _977;
    assign _983 = ~ _982;
    assign _978 = 65'b00000000000000001101101110111000110010110111111000101000000111100;
    assign _977 = { gnd,
                    _10 };
    assign _979 = _977 < _978;
    assign _980 = ~ _979;
    assign _984 = _980 & _983;
    assign _972 = 65'b00000000000000001100100011011110010011001100100111000000101100101;
    assign _973 = _972 < _968;
    assign _974 = ~ _973;
    assign _969 = 65'b00000000000000001100010100010101110100111010000111111110100101101;
    assign _968 = { gnd,
                    _10 };
    assign _970 = _968 < _969;
    assign _971 = ~ _970;
    assign _975 = _971 & _974;
    assign _963 = 65'b00000000000000001101111001000000110001001110000100011111110101000;
    assign _964 = _963 < _959;
    assign _965 = ~ _964;
    assign _960 = 65'b00000000000000001101111000010111011111001001010011110101111111101;
    assign _959 = { gnd,
                    _10 };
    assign _961 = _959 < _960;
    assign _962 = ~ _961;
    assign _966 = _962 & _965;
    assign _954 = 65'b00000000000000001110001010011110010110010110110011111101110101111;
    assign _955 = _954 < _950;
    assign _956 = ~ _955;
    assign _951 = 65'b00000000000000001110000011111110000111111001010010101010100000000;
    assign _950 = { gnd,
                    _10 };
    assign _952 = _950 < _951;
    assign _953 = ~ _952;
    assign _957 = _953 & _956;
    assign _945 = 65'b00000000000000000011000010011011011000111010111001100011110011111;
    assign _946 = _945 < _941;
    assign _947 = ~ _946;
    assign _941 = { gnd,
                    _10 };
    assign _943 = _941 < _1386;
    assign _944 = ~ _943;
    assign _948 = _944 & _947;
    assign _936 = 65'b00000000000000001100011100110101111001001100101110100100111111010;
    assign _937 = _936 < _932;
    assign _938 = ~ _937;
    assign _933 = 65'b00000000000000001100010111011000101101010011010101000111100010111;
    assign _932 = { gnd,
                    _10 };
    assign _934 = _932 < _933;
    assign _935 = ~ _934;
    assign _939 = _935 & _938;
    assign _927 = 65'b00000000000000000010111110111101000111000010010110111001011101110;
    assign _928 = _927 < _923;
    assign _929 = ~ _928;
    assign _924 = 65'b00000000000000000010111101100110111111001111011101110110110111110;
    assign _923 = { gnd,
                    _10 };
    assign _925 = _923 < _924;
    assign _926 = ~ _925;
    assign _930 = _926 & _929;
    assign _918 = 65'b00000000000000000011111110100010100100111111000111101100100010100;
    assign _919 = _918 < _914;
    assign _920 = ~ _919;
    assign _914 = { gnd,
                    _10 };
    assign _916 = _914 < _918;
    assign _917 = ~ _916;
    assign _921 = _917 & _920;
    assign _909 = 65'b00000000000000001000001111101110101111001011101010100100001111100;
    assign _910 = _909 < _905;
    assign _911 = ~ _910;
    assign _906 = 65'b00000000000000001000001000000111110111111000011110011100111100110;
    assign _905 = { gnd,
                    _10 };
    assign _907 = _905 < _906;
    assign _908 = ~ _907;
    assign _912 = _908 & _911;
    assign _900 = 65'b00000000000000000001101000001010011010011000001101111101111101101;
    assign _901 = _900 < _896;
    assign _902 = ~ _901;
    assign _897 = 65'b00000000000000000001011111001011000100011010001101111110110110100;
    assign _896 = { gnd,
                    _10 };
    assign _898 = _896 < _897;
    assign _899 = ~ _898;
    assign _903 = _899 & _902;
    assign _891 = 65'b00000000000000001101100101000000010001110100111110100100011101010;
    assign _892 = _891 < _887;
    assign _893 = ~ _892;
    assign _888 = 65'b00000000000000001101100010101001100001000001100010100001101101111;
    assign _887 = { gnd,
                    _10 };
    assign _889 = _887 < _888;
    assign _890 = ~ _889;
    assign _894 = _890 & _893;
    assign _882 = 65'b00000000000000001011111001100010001010011001010101110001011001100;
    assign _883 = _882 < _878;
    assign _884 = ~ _883;
    assign _879 = 65'b00000000000000001011110101100001101100011100011101011000000010011;
    assign _878 = { gnd,
                    _10 };
    assign _880 = _878 < _879;
    assign _881 = ~ _880;
    assign _885 = _881 & _884;
    assign _873 = 65'b00000000000000001001010111100010100000000001111010101010011111111;
    assign _874 = _873 < _869;
    assign _875 = ~ _874;
    assign _870 = 65'b00000000000000001001010111001010010111010000000011011001100100010;
    assign _869 = { gnd,
                    _10 };
    assign _871 = _869 < _870;
    assign _872 = ~ _871;
    assign _876 = _872 & _875;
    assign _864 = 65'b00000000000000001001001100001010110100010011000010110111000001111;
    assign _865 = _864 < _860;
    assign _866 = ~ _865;
    assign _861 = 65'b00000000000000001001001010101111010000100010010000001101111000000;
    assign _860 = { gnd,
                    _10 };
    assign _862 = _860 < _861;
    assign _863 = ~ _862;
    assign _867 = _863 & _866;
    assign _856 = _1413 < _851;
    assign _857 = ~ _856;
    assign _852 = 65'b00000000000000001011100010001000101011000000100100110000010001100;
    assign _851 = { gnd,
                    _10 };
    assign _853 = _851 < _852;
    assign _854 = ~ _853;
    assign _858 = _854 & _857;
    assign _846 = 65'b00000000000000000100100000110111101000001001011111010101110010111;
    assign _847 = _846 < _842;
    assign _848 = ~ _847;
    assign _843 = 65'b00000000000000000100011110001001001100001111001000011111001111100;
    assign _842 = { gnd,
                    _10 };
    assign _844 = _842 < _843;
    assign _845 = ~ _844;
    assign _849 = _845 & _848;
    assign _837 = 65'b00000000000000000011001101111000011001111101001000110100100110000;
    assign _838 = _837 < _833;
    assign _839 = ~ _838;
    assign _833 = { gnd,
                    _10 };
    assign _835 = _833 < _837;
    assign _836 = ~ _835;
    assign _840 = _836 & _839;
    assign _829 = _945 < _824;
    assign _830 = ~ _829;
    assign _824 = { gnd,
                    _10 };
    assign _826 = _824 < _1383;
    assign _827 = ~ _826;
    assign _831 = _827 & _830;
    assign _819 = 65'b00000000000000000110111110001000100101101000101101111101000111111;
    assign _820 = _819 < _815;
    assign _821 = ~ _820;
    assign _816 = 65'b00000000000000000110110111101101101100110000100011101111111101101;
    assign _815 = { gnd,
                    _10 };
    assign _817 = _815 < _816;
    assign _818 = ~ _817;
    assign _822 = _818 & _821;
    assign _810 = 65'b00000000000000001000110010010111101111111011001001100010110110100;
    assign _811 = _810 < _806;
    assign _812 = ~ _811;
    assign _807 = 65'b00000000000000001000101111001101111010100011001110010100011000110;
    assign _806 = { gnd,
                    _10 };
    assign _808 = _806 < _807;
    assign _809 = ~ _808;
    assign _813 = _809 & _812;
    assign _801 = 65'b00000000000000000100011011110111110000010110100001001100110010000;
    assign _802 = _801 < _797;
    assign _803 = ~ _802;
    assign _798 = 65'b00000000000000000100011001001011110111011110000101101000011000001;
    assign _797 = { gnd,
                    _10 };
    assign _799 = _797 < _798;
    assign _800 = ~ _799;
    assign _804 = _800 & _803;
    assign _792 = 65'b00000000000000001101011010001110000100001111111000000011100011011;
    assign _793 = _792 < _788;
    assign _794 = ~ _793;
    assign _789 = 65'b00000000000000001101010010011001010011110000010010001110000111010;
    assign _788 = { gnd,
                    _10 };
    assign _790 = _788 < _789;
    assign _791 = ~ _790;
    assign _795 = _791 & _794;
    assign _784 = _1278 < _779;
    assign _785 = ~ _784;
    assign _780 = 65'b00000000000000001000111111101100110010010010100011100001011111110;
    assign _779 = { gnd,
                    _10 };
    assign _781 = _779 < _780;
    assign _782 = ~ _781;
    assign _786 = _782 & _785;
    assign _774 = 65'b00000000000000001001010000110001111100000110101011101000111110110;
    assign _775 = _774 < _770;
    assign _776 = ~ _775;
    assign _771 = 65'b00000000000000001001001111001001000011110110011010110110100010100;
    assign _770 = { gnd,
                    _10 };
    assign _772 = _770 < _771;
    assign _773 = ~ _772;
    assign _777 = _773 & _776;
    assign _766 = _1251 < _761;
    assign _767 = ~ _766;
    assign _762 = 65'b00000000000000001101111110100000100010001101000111111111111000101;
    assign _761 = { gnd,
                    _10 };
    assign _763 = _761 < _762;
    assign _764 = ~ _763;
    assign _768 = _764 & _767;
    assign _756 = 65'b00000000000000000000001100111111000110000011011101011111101100000;
    assign _757 = _756 < _752;
    assign _758 = ~ _757;
    assign _753 = 65'b00000000000000000000001011010001111001101001011001011001010000110;
    assign _752 = { gnd,
                    _10 };
    assign _754 = _752 < _753;
    assign _755 = ~ _754;
    assign _759 = _755 & _758;
    assign _747 = 65'b00000000000000000000001011010001111001101001011001011001010000101;
    assign _748 = _747 < _743;
    assign _749 = ~ _748;
    assign _744 = 65'b00000000000000000000000000111010101010110000010100111110100001100;
    assign _743 = { gnd,
                    _10 };
    assign _745 = _743 < _744;
    assign _746 = ~ _745;
    assign _750 = _746 & _749;
    assign _738 = 65'b00000000000000000111011001000100110001110101000110001110010001001;
    assign _739 = _738 < _734;
    assign _740 = ~ _739;
    assign _735 = 65'b00000000000000000111001010101111001011000010001111000001011111000;
    assign _734 = { gnd,
                    _10 };
    assign _736 = _734 < _735;
    assign _737 = ~ _736;
    assign _741 = _737 & _740;
    assign _729 = 65'b00000000000000001010000010000010111001011101101101111100010110000;
    assign _730 = _729 < _725;
    assign _731 = ~ _730;
    assign _725 = { gnd,
                    _10 };
    assign _727 = _725 < _729;
    assign _728 = ~ _727;
    assign _732 = _728 & _731;
    assign _720 = 65'b00000000000000001101100110101011010000111111110001111000101011101;
    assign _721 = _720 < _716;
    assign _722 = ~ _721;
    assign _717 = 65'b00000000000000001101100100010110101010000111100110000000001111001;
    assign _716 = { gnd,
                    _10 };
    assign _718 = _716 < _717;
    assign _719 = ~ _718;
    assign _723 = _719 & _722;
    assign _711 = 65'b00000000000000001111000100101010011100001001000011110100001101010;
    assign _712 = _711 < _707;
    assign _713 = ~ _712;
    assign _708 = 65'b00000000000000001110111101000010101001000100010101100100010000001;
    assign _707 = { gnd,
                    _10 };
    assign _709 = _707 < _708;
    assign _710 = ~ _709;
    assign _714 = _710 & _713;
    assign _702 = 65'b00000000000000000010111100100101111001000110010111111110011011111;
    assign _703 = _702 < _698;
    assign _704 = ~ _703;
    assign _698 = { gnd,
                    _10 };
    assign _700 = _698 < _1323;
    assign _701 = ~ _700;
    assign _705 = _701 & _704;
    assign _693 = 65'b00000000000000001101101010010010000010001101001001001100111100101;
    assign _694 = _693 < _689;
    assign _695 = ~ _694;
    assign _690 = 65'b00000000000000001101100111100111101101110110000111110001011100111;
    assign _689 = { gnd,
                    _10 };
    assign _691 = _689 < _690;
    assign _692 = ~ _691;
    assign _696 = _692 & _695;
    assign _684 = 65'b00000000000000000001111110111001100110001000110111110110001101100;
    assign _685 = _684 < _680;
    assign _686 = ~ _685;
    assign _681 = 65'b00000000000000000001110001010001000000110111101101001111111000100;
    assign _680 = { gnd,
                    _10 };
    assign _682 = _680 < _681;
    assign _683 = ~ _682;
    assign _687 = _683 & _686;
    assign _675 = 65'b00000000000000000000111101100001011000111100001111010100010111100;
    assign _676 = _675 < _671;
    assign _677 = ~ _676;
    assign _672 = 65'b00000000000000000000111010111011101000101100111100001011001111101;
    assign _671 = { gnd,
                    _10 };
    assign _673 = _671 < _672;
    assign _674 = ~ _673;
    assign _678 = _674 & _677;
    assign _666 = 65'b00000000000000001001111100000001100100101001011010000111011110010;
    assign _667 = _666 < _662;
    assign _668 = ~ _667;
    assign _662 = { gnd,
                    _10 };
    assign _664 = _662 < _1104;
    assign _665 = ~ _664;
    assign _669 = _665 & _668;
    assign _657 = 65'b00000000000000000100111001111111100010001011111100010101100011100;
    assign _658 = _657 < _653;
    assign _659 = ~ _658;
    assign _653 = { gnd,
                    _10 };
    assign _655 = _653 < _1527;
    assign _656 = ~ _655;
    assign _660 = _656 & _659;
    assign _648 = 65'b00000000000000001001011110001110011001000111011110101111110110011;
    assign _649 = _648 < _644;
    assign _650 = ~ _649;
    assign _645 = 65'b00000000000000001001011100000010001110100100100000010000111100011;
    assign _644 = { gnd,
                    _10 };
    assign _646 = _644 < _645;
    assign _647 = ~ _646;
    assign _651 = _647 & _650;
    assign _639 = 65'b00000000000000000110001110111111100000101110001100011101100110010;
    assign _640 = _639 < _635;
    assign _641 = ~ _640;
    assign _636 = 65'b00000000000000000110001000101011100111100100000000111110000110100;
    assign _635 = { gnd,
                    _10 };
    assign _637 = _635 < _636;
    assign _638 = ~ _637;
    assign _642 = _638 & _641;
    assign _630 = 65'b00000000000000001110001111000111100001110011000111000101101111100;
    assign _631 = _630 < _626;
    assign _632 = ~ _631;
    assign _626 = { gnd,
                    _10 };
    assign _628 = _626 < _951;
    assign _629 = ~ _628;
    assign _633 = _629 & _632;
    assign _621 = 65'b00000000000000000010111010000111000110100111111000011101110011011;
    assign _622 = _621 < _617;
    assign _623 = ~ _622;
    assign _618 = 65'b00000000000000000010111000110000100001111110010011011001100011110;
    assign _617 = { gnd,
                    _10 };
    assign _619 = _617 < _618;
    assign _620 = ~ _619;
    assign _624 = _620 & _623;
    assign _612 = 65'b00000000000000000001000111001000100001111000000111011011011100000;
    assign _613 = _612 < _608;
    assign _614 = ~ _613;
    assign _609 = 65'b00000000000000000001000100000100101111111110000110101010111010001;
    assign _608 = { gnd,
                    _10 };
    assign _610 = _608 < _609;
    assign _611 = ~ _610;
    assign _615 = _611 & _614;
    assign _604 = _1401 < _599;
    assign _605 = ~ _604;
    assign _599 = { gnd,
                    _10 };
    assign _601 = _599 < _1401;
    assign _602 = ~ _601;
    assign _606 = _602 & _605;
    assign _595 = _1359 < _590;
    assign _596 = ~ _595;
    assign _591 = 65'b00000000000000000100110111010000101010010100010100001001111111011;
    assign _590 = { gnd,
                    _10 };
    assign _592 = _590 < _591;
    assign _593 = ~ _592;
    assign _597 = _593 & _596;
    assign _585 = 65'b00000000000000000101000011101110000101000001010111010100001011010;
    assign _586 = _585 < _581;
    assign _587 = ~ _586;
    assign _582 = 65'b00000000000000000101000011010110111100101010001111101010111110110;
    assign _581 = { gnd,
                    _10 };
    assign _583 = _581 < _582;
    assign _584 = ~ _583;
    assign _588 = _584 & _587;
    assign _576 = 65'b00000000000000000100110100111011111111000101111011000101010001110;
    assign _577 = _576 < _572;
    assign _578 = ~ _577;
    assign _573 = 65'b00000000000000000100101010011101000000101101011000101110111101111;
    assign _572 = { gnd,
                    _10 };
    assign _574 = _572 < _573;
    assign _575 = ~ _574;
    assign _579 = _575 & _578;
    assign _567 = 65'b00000000000000001101011110001100111010011101101011001110000100011;
    assign _568 = _567 < _563;
    assign _569 = ~ _568;
    assign _564 = 65'b00000000000000001101011011101011110010110111110101000011001100100;
    assign _563 = { gnd,
                    _10 };
    assign _565 = _563 < _564;
    assign _566 = ~ _565;
    assign _570 = _566 & _569;
    assign _559 = _1626 < _554;
    assign _560 = ~ _559;
    assign _554 = { gnd,
                    _10 };
    assign _556 = _554 < _1626;
    assign _557 = ~ _556;
    assign _561 = _557 & _560;
    assign _549 = 65'b00000000000000000001010011100000001101010001010001100110011100011;
    assign _550 = _549 < _545;
    assign _551 = ~ _550;
    assign _546 = 65'b00000000000000000001001100001010111001001110100110011000001000010;
    assign _545 = { gnd,
                    _10 };
    assign _547 = _545 < _546;
    assign _548 = ~ _547;
    assign _552 = _548 & _551;
    assign _541 = _1608 < _536;
    assign _542 = ~ _541;
    assign _536 = { gnd,
                    _10 };
    assign _538 = _536 < _1608;
    assign _539 = ~ _538;
    assign _543 = _539 & _542;
    assign _532 = _1059 < _527;
    assign _533 = ~ _532;
    assign _528 = 65'b00000000000000001001001001111001100100011001011000111100101110110;
    assign _527 = { gnd,
                    _10 };
    assign _529 = _527 < _528;
    assign _530 = ~ _529;
    assign _534 = _530 & _533;
    assign _522 = 65'b00000000000000000101010011100010111110010101001101011111001111100;
    assign _523 = _522 < _518;
    assign _524 = ~ _523;
    assign _519 = 65'b00000000000000000101010000000111001000011101001011011001101011000;
    assign _518 = { gnd,
                    _10 };
    assign _520 = _518 < _519;
    assign _521 = ~ _520;
    assign _525 = _521 & _524;
    assign _513 = 65'b00000000000000000101111101101111111000000101010100110110111011001;
    assign _514 = _513 < _509;
    assign _515 = ~ _514;
    assign _510 = 65'b00000000000000000101110101010111100010101101011010010111010000111;
    assign _509 = { gnd,
                    _10 };
    assign _511 = _509 < _510;
    assign _512 = ~ _511;
    assign _516 = _512 & _515;
    assign _505 = _1494 < _500;
    assign _506 = ~ _505;
    assign _500 = { gnd,
                    _10 };
    assign _502 = _500 < _1491;
    assign _503 = ~ _502;
    assign _507 = _503 & _506;
    assign _495 = 65'b00000000000000000100111010011101100101101111100010110110001111011;
    assign _496 = _495 < _491;
    assign _497 = ~ _496;
    assign _491 = { gnd,
                    _10 };
    assign _493 = _491 < _657;
    assign _494 = ~ _493;
    assign _498 = _494 & _497;
    assign _487 = _639 < _482;
    assign _488 = ~ _487;
    assign _483 = 65'b00000000000000000110000100100101001010111100011110011000000010111;
    assign _482 = { gnd,
                    _10 };
    assign _484 = _482 < _483;
    assign _485 = ~ _484;
    assign _489 = _485 & _488;
    assign _477 = 65'b00000000000000000001011000001100011010001111100011010001001100101;
    assign _478 = _477 < _473;
    assign _479 = ~ _478;
    assign _474 = 65'b00000000000000000001010000000111001011101000011011001111001010001;
    assign _473 = { gnd,
                    _10 };
    assign _475 = _473 < _474;
    assign _476 = ~ _475;
    assign _480 = _476 & _479;
    assign _468 = 65'b00000000000000001111010011101000011110100100100100010011110100110;
    assign _469 = _468 < _464;
    assign _470 = ~ _469;
    assign _465 = 65'b00000000000000001111001101001010011110011100110010111010000000011;
    assign _464 = { gnd,
                    _10 };
    assign _466 = _464 < _465;
    assign _467 = ~ _466;
    assign _471 = _467 & _470;
    assign _459 = 65'b00000000000000000101001000011011001110000111111010110100011101011;
    assign _460 = _459 < _455;
    assign _461 = ~ _460;
    assign _456 = 65'b00000000000000000101000111010111110100000011010010011101010111101;
    assign _455 = { gnd,
                    _10 };
    assign _457 = _455 < _456;
    assign _458 = ~ _457;
    assign _462 = _458 & _461;
    assign _450 = 65'b00000000000000001000101111001101111010100011001110010100011000101;
    assign _451 = _450 < _446;
    assign _452 = ~ _451;
    assign _447 = 65'b00000000000000001000100101111101110001010111100010101110001001111;
    assign _446 = { gnd,
                    _10 };
    assign _448 = _446 < _447;
    assign _449 = ~ _448;
    assign _453 = _449 & _452;
    assign _442 = _459 < _437;
    assign _443 = ~ _442;
    assign _437 = { gnd,
                    _10 };
    assign _439 = _437 < _1593;
    assign _440 = ~ _439;
    assign _444 = _440 & _443;
    assign _432 = 65'b00000000000000001101111100111010100011000101101011111100100101000;
    assign _433 = _432 < _428;
    assign _434 = ~ _433;
    assign _429 = 65'b00000000000000001101111100100010000010010100101101000010110001001;
    assign _428 = { gnd,
                    _10 };
    assign _430 = _428 < _429;
    assign _431 = ~ _430;
    assign _435 = _431 & _434;
    assign _424 = _918 < _419;
    assign _425 = ~ _424;
    assign _420 = 65'b00000000000000000011110010101100101101111101011100010000111111000;
    assign _419 = { gnd,
                    _10 };
    assign _421 = _419 < _420;
    assign _422 = ~ _421;
    assign _426 = _422 & _425;
    assign _415 = _576 < _410;
    assign _416 = ~ _415;
    assign _410 = { gnd,
                    _10 };
    assign _412 = _410 < _573;
    assign _413 = ~ _412;
    assign _417 = _413 & _416;
    assign _405 = 65'b00000000000000000001000011001001101000010011101001001010110111100;
    assign _406 = _405 < _401;
    assign _407 = ~ _406;
    assign _402 = 65'b00000000000000000001000000011010010011001000000100010111001010000;
    assign _401 = { gnd,
                    _10 };
    assign _403 = _401 < _402;
    assign _404 = ~ _403;
    assign _408 = _404 & _407;
    assign _396 = 65'b00000000000000001110111101000010101001000100010101100100010000000;
    assign _397 = _396 < _392;
    assign _398 = ~ _397;
    assign _392 = { gnd,
                    _10 };
    assign _394 = _392 < _396;
    assign _395 = ~ _394;
    assign _399 = _395 & _398;
    assign _387 = 65'b00000000000000000100111111101001111111111000100100011010001001100;
    assign _388 = _387 < _383;
    assign _389 = ~ _388;
    assign _384 = 65'b00000000000000000100111111000010010111001100101011010011011100010;
    assign _383 = { gnd,
                    _10 };
    assign _385 = _383 < _384;
    assign _386 = ~ _385;
    assign _390 = _386 & _389;
    assign _378 = 65'b00000000000000000011000011100110111001001100110111011110100000001;
    assign _379 = _378 < _374;
    assign _380 = ~ _379;
    assign _374 = { gnd,
                    _10 };
    assign _376 = _374 < _945;
    assign _377 = ~ _376;
    assign _381 = _377 & _380;
    assign _369 = 65'b00000000000000001110110101001001111110110101101110010001000011111;
    assign _370 = _369 < _365;
    assign _371 = ~ _370;
    assign _366 = 65'b00000000000000001110100101100101110111001100010010110101010101001;
    assign _365 = { gnd,
                    _10 };
    assign _367 = _365 < _366;
    assign _368 = ~ _367;
    assign _372 = _368 & _371;
    assign _360 = 65'b00000000000000001101100001011111110101100011101111111101111110101;
    assign _361 = _360 < _356;
    assign _362 = ~ _361;
    assign _357 = 65'b00000000000000001101011111011010100010000111010111100000101110110;
    assign _356 = { gnd,
                    _10 };
    assign _358 = _356 < _357;
    assign _359 = ~ _358;
    assign _363 = _359 & _362;
    assign _351 = 65'b00000000000000000101000111110101011000001010110001111100110001100;
    assign _352 = _351 < _347;
    assign _353 = ~ _352;
    assign _348 = 65'b00000000000000000101000110100100110001000110001100000100101000111;
    assign _347 = { gnd,
                    _10 };
    assign _349 = _347 < _348;
    assign _350 = ~ _349;
    assign _354 = _350 & _353;
    assign _342 = 65'b00000000000000001001101010000100100111100000010001111000001010101;
    assign _343 = _342 < _338;
    assign _344 = ~ _343;
    assign _339 = 65'b00000000000000001001100111010001001001100111111100101011110010100;
    assign _338 = { gnd,
                    _10 };
    assign _340 = _338 < _339;
    assign _341 = ~ _340;
    assign _345 = _341 & _344;
    assign _333 = 65'b00000000000000000100011111011110010011101100101100100101101110011;
    assign _334 = _333 < _329;
    assign _335 = ~ _334;
    assign _330 = 65'b00000000000000000100011100111110010001000001001010001001101010111;
    assign _329 = { gnd,
                    _10 };
    assign _331 = _329 < _330;
    assign _332 = ~ _331;
    assign _336 = _332 & _335;
    assign _325 = _927 < _320;
    assign _326 = ~ _325;
    assign _320 = { gnd,
                    _10 };
    assign _322 = _320 < _924;
    assign _323 = ~ _322;
    assign _327 = _323 & _326;
    assign _315 = 65'b00000000000000001000001100001001100001111111010111001111010011111;
    assign _316 = _315 < _311;
    assign _317 = ~ _316;
    assign _312 = 65'b00000000000000001000000011000000000000110111001100000111001100000;
    assign _311 = { gnd,
                    _10 };
    assign _313 = _311 < _312;
    assign _314 = ~ _313;
    assign _318 = _314 & _317;
    assign _307 = _1590 < _302;
    assign _308 = ~ _307;
    assign _303 = 65'b00000000000000000101000101001010101000110100010111101010000011011;
    assign _302 = { gnd,
                    _10 };
    assign _304 = _302 < _303;
    assign _305 = ~ _304;
    assign _309 = _305 & _308;
    assign _297 = 65'b00000000000000000000110101010111001011110001010101110001110110001;
    assign _298 = _297 < _293;
    assign _299 = ~ _298;
    assign _294 = 65'b00000000000000000000100110010000011000111011100001001000100000111;
    assign _293 = { gnd,
                    _10 };
    assign _295 = _293 < _294;
    assign _296 = ~ _295;
    assign _300 = _296 & _299;
    assign _288 = 65'b00000000000000001001001110110010010001001000101111100000010101111;
    assign _289 = _288 < _284;
    assign _290 = ~ _289;
    assign _285 = 65'b00000000000000001001001110000000000000010000100100001001010000010;
    assign _284 = { gnd,
                    _10 };
    assign _286 = _284 < _285;
    assign _287 = ~ _286;
    assign _291 = _287 & _290;
    assign _279 = 65'b00000000000000001011111110101011000000111111011100101110110111111;
    assign _280 = _279 < _275;
    assign _281 = ~ _280;
    assign _276 = 65'b00000000000000001011101111011101001000001100010001010100000110100;
    assign _275 = { gnd,
                    _10 };
    assign _277 = _275 < _276;
    assign _278 = ~ _277;
    assign _282 = _278 & _281;
    assign _270 = 65'b00000000000000001001101000000101110100011011011111110011010011001;
    assign _271 = _270 < _266;
    assign _272 = ~ _271;
    assign _267 = 65'b00000000000000001001100101111100001111011000100110010100101110100;
    assign _266 = { gnd,
                    _10 };
    assign _268 = _266 < _267;
    assign _269 = ~ _268;
    assign _273 = _269 & _272;
    assign _262 = _1260 < _257;
    assign _263 = ~ _262;
    assign _258 = 65'b00000000000000001100000101011110101111111001111000001000010110001;
    assign _257 = { gnd,
                    _10 };
    assign _259 = _257 < _258;
    assign _260 = ~ _259;
    assign _264 = _260 & _263;
    assign _253 = _582 < _248;
    assign _254 = ~ _253;
    assign _249 = 65'b00000000000000000101000011000111101110100010010010100110110110110;
    assign _248 = { gnd,
                    _10 };
    assign _250 = _248 < _249;
    assign _251 = ~ _250;
    assign _255 = _251 & _254;
    assign _243 = 65'b00000000000000001010001110101010010010010100101011000010001100001;
    assign _244 = _243 < _239;
    assign _245 = ~ _244;
    assign _239 = { gnd,
                    _10 };
    assign _241 = _239 < _729;
    assign _242 = ~ _241;
    assign _246 = _242 & _245;
    assign _234 = 65'b00000000000000000100100010010100001101110011100110100110110000110;
    assign _235 = _234 < _230;
    assign _236 = ~ _235;
    assign _231 = 65'b00000000000000000100100000000010110101100100011011000010110001100;
    assign _230 = { gnd,
                    _10 };
    assign _232 = _230 < _231;
    assign _233 = ~ _232;
    assign _237 = _233 & _236;
    assign _226 = _684 < _221;
    assign _227 = ~ _226;
    assign _222 = 65'b00000000000000000001111000010000000000101110000100111010100011101;
    assign _221 = { gnd,
                    _10 };
    assign _223 = _221 < _222;
    assign _224 = ~ _223;
    assign _228 = _224 & _227;
    assign _216 = 65'b00000000000000000111000011111010010011011101010001111101001000011;
    assign _217 = _216 < _212;
    assign _218 = ~ _217;
    assign _213 = 65'b00000000000000000110111110001000100101101000101101111101001000000;
    assign _212 = { gnd,
                    _10 };
    assign _214 = _212 < _213;
    assign _215 = ~ _214;
    assign _219 = _215 & _218;
    assign _208 = _963 < _203;
    assign _209 = ~ _208;
    assign _203 = { gnd,
                    _10 };
    assign _205 = _203 < _960;
    assign _206 = ~ _205;
    assign _210 = _206 & _209;
    assign _198 = 65'b00000000000000000010010000011001100000100000110110111111000000001;
    assign _199 = _198 < _194;
    assign _200 = ~ _199;
    assign _194 = { gnd,
                    _10 };
    assign _196 = _194 < _1329;
    assign _197 = ~ _196;
    assign _201 = _197 & _200;
    assign _189 = 65'b00000000000000000000111011111101100010100101100101111000011000100;
    assign _190 = _189 < _185;
    assign _191 = ~ _190;
    assign _186 = 65'b00000000000000000000111000111000001100010011010111111011010110100;
    assign _185 = { gnd,
                    _10 };
    assign _187 = _185 < _186;
    assign _188 = ~ _187;
    assign _192 = _188 & _191;
    assign _180 = 65'b00000000000000001110100001010111110111110100010110101100000100101;
    assign _181 = _180 < _176;
    assign _182 = ~ _181;
    assign _177 = 65'b00000000000000001110011010010110000101010111001000110000000011010;
    assign _176 = { gnd,
                    _10 };
    assign _178 = _176 < _177;
    assign _179 = ~ _178;
    assign _183 = _179 & _182;
    assign _172 = _1503 < _167;
    assign _173 = ~ _172;
    assign _167 = { gnd,
                    _10 };
    assign _169 = _167 < _1500;
    assign _170 = ~ _169;
    assign _174 = _170 & _173;
    assign _162 = 65'b00000000000000001101101011100111100111100100100111010101110110010;
    assign _163 = _162 < _158;
    assign _164 = ~ _163;
    assign _159 = 65'b00000000000000001101101001011100011101100111000010010010010100000;
    assign _158 = { gnd,
                    _10 };
    assign _160 = _158 < _159;
    assign _161 = ~ _160;
    assign _165 = _161 & _164;
    assign _153 = 65'b00000000000000000011000001100000100011000111001010101000101100000;
    assign _154 = _153 < _149;
    assign _155 = ~ _154;
    assign _150 = 65'b00000000000000000011000000010100010011110010101111010110110011110;
    assign _149 = { gnd,
                    _10 };
    assign _151 = _149 < _150;
    assign _152 = ~ _151;
    assign _156 = _152 & _155;
    assign _145 = _150 < _140;
    assign _146 = ~ _145;
    assign _140 = { gnd,
                    _10 };
    assign _142 = _140 < _927;
    assign _143 = ~ _142;
    assign _147 = _143 & _146;
    assign _135 = 65'b00000000000000000000111111010001000011000001100100000010111111010;
    assign _136 = _135 < _131;
    assign _137 = ~ _136;
    assign _132 = 65'b00000000000000000000111100011100010101111001101011011110001100000;
    assign _131 = { gnd,
                    _10 };
    assign _133 = _131 < _132;
    assign _134 = ~ _133;
    assign _138 = _134 & _137;
    assign _126 = 65'b00000000000000001001011010000000010111100000100000111010100001110;
    assign _127 = _126 < _122;
    assign _128 = ~ _127;
    assign _122 = { gnd,
                    _10 };
    assign _124 = _122 < _1482;
    assign _125 = ~ _124;
    assign _129 = _125 & _128;
    assign _118 = _369 < _113;
    assign _119 = ~ _118;
    assign _113 = { gnd,
                    _10 };
    assign _115 = _113 < _366;
    assign _116 = ~ _115;
    assign _120 = _116 & _119;
    assign _108 = 65'b00000000000000000100010000100101010001100101010110000101111111110;
    assign _109 = _108 < _104;
    assign _110 = ~ _109;
    assign _105 = 65'b00000000000000000100000101101010101010000100011000110100101001000;
    assign _104 = { gnd,
                    _10 };
    assign _106 = _104 < _105;
    assign _107 = ~ _106;
    assign _111 = _107 & _110;
    assign _99 = 65'b00000000000000001010011001010000111110010110111101101100000000100;
    assign _100 = _99 < _95;
    assign _101 = ~ _100;
    assign _96 = 65'b00000000000000001010010100011000001011011110001000101101000010001;
    assign _95 = { gnd,
                   _10 };
    assign _97 = _95 < _96;
    assign _98 = ~ _97;
    assign _102 = _98 & _101;
    assign _91 = _378 < _86;
    assign _92 = ~ _91;
    assign _86 = { gnd,
                   _10 };
    assign _88 = _86 < _1386;
    assign _89 = ~ _88;
    assign _93 = _89 & _92;
    assign _81 = 65'b00000000000000001001100011010001001100110000110110001100011110000;
    assign _82 = _81 < _77;
    assign _83 = ~ _82;
    assign _78 = 65'b00000000000000001001100000100100100001110101110101010101010110010;
    assign _77 = { gnd,
                   _10 };
    assign _79 = _77 < _78;
    assign _80 = ~ _79;
    assign _84 = _80 & _83;
    assign _72 = 65'b00000000000000000100011000110001111001100110100000100011110111110;
    assign _73 = _72 < _68;
    assign _74 = ~ _73;
    assign _69 = 65'b00000000000000000100010110000100001111000000101010111010100111011;
    assign _68 = { gnd,
                   _10 };
    assign _70 = _68 < _69;
    assign _71 = ~ _70;
    assign _75 = _71 & _74;
    assign _63 = 65'b00000000000000000111101111111110001101101101110010001101100011010;
    assign _64 = _63 < _59;
    assign _65 = ~ _64;
    assign _59 = { gnd,
                   _10 };
    assign _61 = _59 < _63;
    assign _62 = ~ _61;
    assign _66 = _62 & _65;
    assign _55 = _1599 < _50;
    assign _56 = ~ _55;
    assign _50 = { gnd,
                   _10 };
    assign _52 = _50 < _1440;
    assign _53 = ~ _52;
    assign _57 = _53 & _56;
    assign _46 = _285 < _41;
    assign _47 = ~ _46;
    assign _42 = 65'b00000000000000001001001101101000011011110101010000010111001101100;
    assign _41 = { gnd,
                   _10 };
    assign _43 = _41 < _42;
    assign _44 = ~ _43;
    assign _48 = _44 & _47;
    assign _36 = 65'b00000000000000001111011000001000000111000100101001100000010001011;
    assign _37 = _36 < _32;
    assign _38 = ~ _37;
    assign _33 = 65'b00000000000000001111010001001010001100100001001101101001111011000;
    assign _32 = { gnd,
                   _10 };
    assign _34 = _32 < _33;
    assign _35 = ~ _34;
    assign _39 = _35 & _38;
    assign _28 = _1125 < _23;
    assign _29 = ~ _28;
    assign _24 = 65'b00000000000000001001010011111100110010010010111001011111011001111;
    assign _23 = { gnd,
                   _10 };
    assign _25 = _23 < _24;
    assign _26 = ~ _25;
    assign _30 = _26 & _29;
    assign _19 = 65'b00000000000000001101110001010100101000010000100110011000010000000;
    assign _20 = _19 < _15;
    assign _21 = ~ _20;
    assign _16 = 65'b00000000000000001101110000101011000100100001000000100000100000011;
    assign _10 = ingredient_id;
    assign gnd = 1'b0;
    assign _15 = { gnd,
                   _10 };
    assign _17 = _15 < _16;
    assign _18 = ~ _17;
    assign _22 = _18 & _21;
    assign _31 = _22 | _30;
    assign _40 = _31 | _39;
    assign _49 = _40 | _48;
    assign _58 = _49 | _57;
    assign _67 = _58 | _66;
    assign _76 = _67 | _75;
    assign _85 = _76 | _84;
    assign _94 = _85 | _93;
    assign _103 = _94 | _102;
    assign _112 = _103 | _111;
    assign _121 = _112 | _120;
    assign _130 = _121 | _129;
    assign _139 = _130 | _138;
    assign _148 = _139 | _147;
    assign _157 = _148 | _156;
    assign _166 = _157 | _165;
    assign _175 = _166 | _174;
    assign _184 = _175 | _183;
    assign _193 = _184 | _192;
    assign _202 = _193 | _201;
    assign _211 = _202 | _210;
    assign _220 = _211 | _219;
    assign _229 = _220 | _228;
    assign _238 = _229 | _237;
    assign _247 = _238 | _246;
    assign _256 = _247 | _255;
    assign _265 = _256 | _264;
    assign _274 = _265 | _273;
    assign _283 = _274 | _282;
    assign _292 = _283 | _291;
    assign _301 = _292 | _300;
    assign _310 = _301 | _309;
    assign _319 = _310 | _318;
    assign _328 = _319 | _327;
    assign _337 = _328 | _336;
    assign _346 = _337 | _345;
    assign _355 = _346 | _354;
    assign _364 = _355 | _363;
    assign _373 = _364 | _372;
    assign _382 = _373 | _381;
    assign _391 = _382 | _390;
    assign _400 = _391 | _399;
    assign _409 = _400 | _408;
    assign _418 = _409 | _417;
    assign _427 = _418 | _426;
    assign _436 = _427 | _435;
    assign _445 = _436 | _444;
    assign _454 = _445 | _453;
    assign _463 = _454 | _462;
    assign _472 = _463 | _471;
    assign _481 = _472 | _480;
    assign _490 = _481 | _489;
    assign _499 = _490 | _498;
    assign _508 = _499 | _507;
    assign _517 = _508 | _516;
    assign _526 = _517 | _525;
    assign _535 = _526 | _534;
    assign _544 = _535 | _543;
    assign _553 = _544 | _552;
    assign _562 = _553 | _561;
    assign _571 = _562 | _570;
    assign _580 = _571 | _579;
    assign _589 = _580 | _588;
    assign _598 = _589 | _597;
    assign _607 = _598 | _606;
    assign _616 = _607 | _615;
    assign _625 = _616 | _624;
    assign _634 = _625 | _633;
    assign _643 = _634 | _642;
    assign _652 = _643 | _651;
    assign _661 = _652 | _660;
    assign _670 = _661 | _669;
    assign _679 = _670 | _678;
    assign _688 = _679 | _687;
    assign _697 = _688 | _696;
    assign _706 = _697 | _705;
    assign _715 = _706 | _714;
    assign _724 = _715 | _723;
    assign _733 = _724 | _732;
    assign _742 = _733 | _741;
    assign _751 = _742 | _750;
    assign _760 = _751 | _759;
    assign _769 = _760 | _768;
    assign _778 = _769 | _777;
    assign _787 = _778 | _786;
    assign _796 = _787 | _795;
    assign _805 = _796 | _804;
    assign _814 = _805 | _813;
    assign _823 = _814 | _822;
    assign _832 = _823 | _831;
    assign _841 = _832 | _840;
    assign _850 = _841 | _849;
    assign _859 = _850 | _858;
    assign _868 = _859 | _867;
    assign _877 = _868 | _876;
    assign _886 = _877 | _885;
    assign _895 = _886 | _894;
    assign _904 = _895 | _903;
    assign _913 = _904 | _912;
    assign _922 = _913 | _921;
    assign _931 = _922 | _930;
    assign _940 = _931 | _939;
    assign _949 = _940 | _948;
    assign _958 = _949 | _957;
    assign _967 = _958 | _966;
    assign _976 = _967 | _975;
    assign _985 = _976 | _984;
    assign _994 = _985 | _993;
    assign _1003 = _994 | _1002;
    assign _1012 = _1003 | _1011;
    assign _1021 = _1012 | _1020;
    assign _1030 = _1021 | _1029;
    assign _1039 = _1030 | _1038;
    assign _1048 = _1039 | _1047;
    assign _1057 = _1048 | _1056;
    assign _1066 = _1057 | _1065;
    assign _1075 = _1066 | _1074;
    assign _1084 = _1075 | _1083;
    assign _1093 = _1084 | _1092;
    assign _1102 = _1093 | _1101;
    assign _1111 = _1102 | _1110;
    assign _1120 = _1111 | _1119;
    assign _1129 = _1120 | _1128;
    assign _1138 = _1129 | _1137;
    assign _1147 = _1138 | _1146;
    assign _1156 = _1147 | _1155;
    assign _1165 = _1156 | _1164;
    assign _1174 = _1165 | _1173;
    assign _1183 = _1174 | _1182;
    assign _1192 = _1183 | _1191;
    assign _1201 = _1192 | _1200;
    assign _1210 = _1201 | _1209;
    assign _1219 = _1210 | _1218;
    assign _1228 = _1219 | _1227;
    assign _1237 = _1228 | _1236;
    assign _1246 = _1237 | _1245;
    assign _1255 = _1246 | _1254;
    assign _1264 = _1255 | _1263;
    assign _1273 = _1264 | _1272;
    assign _1282 = _1273 | _1281;
    assign _1291 = _1282 | _1290;
    assign _1300 = _1291 | _1299;
    assign _1309 = _1300 | _1308;
    assign _1318 = _1309 | _1317;
    assign _1327 = _1318 | _1326;
    assign _1336 = _1327 | _1335;
    assign _1345 = _1336 | _1344;
    assign _1354 = _1345 | _1353;
    assign _1363 = _1354 | _1362;
    assign _1372 = _1363 | _1371;
    assign _1381 = _1372 | _1380;
    assign _1390 = _1381 | _1389;
    assign _1399 = _1390 | _1398;
    assign _1408 = _1399 | _1407;
    assign _1417 = _1408 | _1416;
    assign _1426 = _1417 | _1425;
    assign _1435 = _1426 | _1434;
    assign _1444 = _1435 | _1443;
    assign _1453 = _1444 | _1452;
    assign _1462 = _1453 | _1461;
    assign _1471 = _1462 | _1470;
    assign _1480 = _1471 | _1479;
    assign _1489 = _1480 | _1488;
    assign _1498 = _1489 | _1497;
    assign _1507 = _1498 | _1506;
    assign _1516 = _1507 | _1515;
    assign _1525 = _1516 | _1524;
    assign _1534 = _1525 | _1533;
    assign _1543 = _1534 | _1542;
    assign _1552 = _1543 | _1551;
    assign _1561 = _1552 | _1560;
    assign _1570 = _1561 | _1569;
    assign _1579 = _1570 | _1578;
    assign _1588 = _1579 | _1587;
    assign _1597 = _1588 | _1596;
    assign _1606 = _1597 | _1605;
    assign _1615 = _1606 | _1614;
    assign _1624 = _1615 | _1623;
    assign _1633 = _1624 | _1632;
    assign _1642 = _1633 | _1641;
    assign _1651 = _1642 | _1650;
    assign _1660 = _1651 | _1659;
    assign _1669 = _1660 | _1668;
    assign _1678 = _1669 | _1677;
    assign _1687 = _1678 | _1686;
    assign _1696 = _1687 | _1695;
    assign is_fresh = _1696;
    assign total_count = _1698;

endmodule
