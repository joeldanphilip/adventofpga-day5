module sorter_and_merger (
    wr_end,
    wr_start,
    wr_enable,
    clear,
    clock,
    start_processing,
    result,
    done_flag,
    state_debug
);

    input [63:0] wr_end;
    input [63:0] wr_start;
    input wr_enable;
    input clear;
    input clock;
    input start_processing;
    output [63:0] result;
    output done_flag;
    output [1:0] state_debug;

    wire _428;
    wire [63:0] _5492;
    wire [63:0] _5495;
    wire _1051;
    wire [63:0] _1052;
    wire [63:0] _1053;
    wire [63:0] _3;
    reg [63:0] _433;
    wire [63:0] _5494;
    wire [63:0] _5496;
    wire [63:0] _5497;
    reg [63:0] _1047;
    wire [64:0] _1048;
    wire [64:0] _5464;
    wire [64:0] _5463;
    wire _5465;
    wire [63:0] _5466;
    wire [63:0] _5;
    wire [63:0] _5457;
    wire [63:0] _4228;
    wire [63:0] _4196;
    wire [63:0] _4164;
    wire [63:0] _4132;
    wire [63:0] _4100;
    wire [63:0] _4068;
    wire [63:0] _4036;
    wire [63:0] _4004;
    wire [63:0] _3972;
    wire [63:0] _3940;
    wire [63:0] _3908;
    wire [63:0] _3876;
    wire [63:0] _3844;
    wire [63:0] _3812;
    wire [63:0] _3780;
    wire [63:0] _3748;
    wire [63:0] _3716;
    wire [63:0] _3684;
    wire [63:0] _3652;
    wire [63:0] _3620;
    wire [63:0] _3588;
    wire [63:0] _3556;
    wire [63:0] _3524;
    wire [63:0] _3492;
    wire [63:0] _3460;
    wire [63:0] _3428;
    wire [63:0] _3396;
    wire [63:0] _3364;
    wire [63:0] _3332;
    wire [63:0] _3300;
    wire [63:0] _3268;
    wire [63:0] _3236;
    wire [63:0] _3204;
    wire [63:0] _3172;
    wire [63:0] _3140;
    wire [63:0] _3108;
    wire [63:0] _3076;
    wire [63:0] _3044;
    wire [63:0] _3012;
    wire [63:0] _2980;
    wire [63:0] _2948;
    wire [63:0] _2916;
    wire [63:0] _2884;
    wire [63:0] _2852;
    wire [63:0] _2820;
    wire [63:0] _2788;
    wire [63:0] _2756;
    wire [63:0] _2724;
    wire [63:0] _2692;
    wire [63:0] _2660;
    wire [63:0] _2628;
    wire [63:0] _2596;
    wire [63:0] _2564;
    wire [63:0] _2532;
    wire [63:0] _2500;
    wire [63:0] _2468;
    wire [63:0] _2436;
    wire [63:0] _2404;
    wire [63:0] _2372;
    wire [63:0] _2340;
    wire [63:0] _2308;
    wire [63:0] _2276;
    wire [63:0] _2244;
    wire [63:0] _2212;
    wire [63:0] _2180;
    wire [63:0] _2148;
    wire [63:0] _2116;
    wire [63:0] _2084;
    wire [63:0] _2052;
    wire [63:0] _2020;
    wire [63:0] _1988;
    wire [63:0] _1956;
    wire [63:0] _1924;
    wire [63:0] _1892;
    wire [63:0] _1860;
    wire [63:0] _1828;
    wire [63:0] _1796;
    wire [63:0] _1764;
    wire [63:0] _1732;
    wire [63:0] _1700;
    wire [63:0] _1668;
    wire [63:0] _1636;
    wire [63:0] _1604;
    wire [63:0] _1572;
    wire [63:0] _1540;
    wire [63:0] _1508;
    wire [63:0] _1476;
    wire [63:0] _1444;
    wire [63:0] _1412;
    wire [63:0] _1380;
    wire [63:0] _1348;
    wire [63:0] _1316;
    wire [63:0] _1284;
    wire [63:0] _1252;
    wire [63:0] _1220;
    wire [63:0] _1188;
    wire [63:0] _1156;
    wire [63:0] _1124;
    wire [63:0] _1092;
    wire [63:0] _1076;
    wire [63:0] _1072;
    wire [63:0] _1077;
    wire [63:0] _1078;
    wire _1056;
    wire [63:0] _1079;
    wire [63:0] _6;
    reg [63:0] _1061;
    wire [63:0] _1085;
    wire [63:0] _1093;
    wire [63:0] _1094;
    wire _1080;
    wire [63:0] _1095;
    wire [63:0] _7;
    reg [63:0] _1071;
    wire [63:0] _1108;
    wire [63:0] _1104;
    wire [63:0] _1109;
    wire [63:0] _1110;
    wire _1096;
    wire [63:0] _1111;
    wire [63:0] _8;
    reg [63:0] _1091;
    wire [63:0] _1117;
    wire [63:0] _1125;
    wire [63:0] _1126;
    wire _1112;
    wire [63:0] _1127;
    wire [63:0] _9;
    reg [63:0] _1103;
    wire [63:0] _1140;
    wire [63:0] _1136;
    wire [63:0] _1141;
    wire [63:0] _1142;
    wire _1128;
    wire [63:0] _1143;
    wire [63:0] _10;
    reg [63:0] _1123;
    wire [63:0] _1149;
    wire [63:0] _1157;
    wire [63:0] _1158;
    wire _1144;
    wire [63:0] _1159;
    wire [63:0] _11;
    reg [63:0] _1135;
    wire [63:0] _1172;
    wire [63:0] _1168;
    wire [63:0] _1173;
    wire [63:0] _1174;
    wire _1160;
    wire [63:0] _1175;
    wire [63:0] _12;
    reg [63:0] _1155;
    wire [63:0] _1181;
    wire [63:0] _1189;
    wire [63:0] _1190;
    wire _1176;
    wire [63:0] _1191;
    wire [63:0] _13;
    reg [63:0] _1167;
    wire [63:0] _1204;
    wire [63:0] _1200;
    wire [63:0] _1205;
    wire [63:0] _1206;
    wire _1192;
    wire [63:0] _1207;
    wire [63:0] _14;
    reg [63:0] _1187;
    wire [63:0] _1213;
    wire [63:0] _1221;
    wire [63:0] _1222;
    wire _1208;
    wire [63:0] _1223;
    wire [63:0] _15;
    reg [63:0] _1199;
    wire [63:0] _1236;
    wire [63:0] _1232;
    wire [63:0] _1237;
    wire [63:0] _1238;
    wire _1224;
    wire [63:0] _1239;
    wire [63:0] _16;
    reg [63:0] _1219;
    wire [63:0] _1245;
    wire [63:0] _1253;
    wire [63:0] _1254;
    wire _1240;
    wire [63:0] _1255;
    wire [63:0] _17;
    reg [63:0] _1231;
    wire [63:0] _1268;
    wire [63:0] _1264;
    wire [63:0] _1269;
    wire [63:0] _1270;
    wire _1256;
    wire [63:0] _1271;
    wire [63:0] _18;
    reg [63:0] _1251;
    wire [63:0] _1277;
    wire [63:0] _1285;
    wire [63:0] _1286;
    wire _1272;
    wire [63:0] _1287;
    wire [63:0] _19;
    reg [63:0] _1263;
    wire [63:0] _1300;
    wire [63:0] _1296;
    wire [63:0] _1301;
    wire [63:0] _1302;
    wire _1288;
    wire [63:0] _1303;
    wire [63:0] _20;
    reg [63:0] _1283;
    wire [63:0] _1309;
    wire [63:0] _1317;
    wire [63:0] _1318;
    wire _1304;
    wire [63:0] _1319;
    wire [63:0] _21;
    reg [63:0] _1295;
    wire [63:0] _1332;
    wire [63:0] _1328;
    wire [63:0] _1333;
    wire [63:0] _1334;
    wire _1320;
    wire [63:0] _1335;
    wire [63:0] _22;
    reg [63:0] _1315;
    wire [63:0] _1341;
    wire [63:0] _1349;
    wire [63:0] _1350;
    wire _1336;
    wire [63:0] _1351;
    wire [63:0] _23;
    reg [63:0] _1327;
    wire [63:0] _1364;
    wire [63:0] _1360;
    wire [63:0] _1365;
    wire [63:0] _1366;
    wire _1352;
    wire [63:0] _1367;
    wire [63:0] _24;
    reg [63:0] _1347;
    wire [63:0] _1373;
    wire [63:0] _1381;
    wire [63:0] _1382;
    wire _1368;
    wire [63:0] _1383;
    wire [63:0] _25;
    reg [63:0] _1359;
    wire [63:0] _1396;
    wire [63:0] _1392;
    wire [63:0] _1397;
    wire [63:0] _1398;
    wire _1384;
    wire [63:0] _1399;
    wire [63:0] _26;
    reg [63:0] _1379;
    wire [63:0] _1405;
    wire [63:0] _1413;
    wire [63:0] _1414;
    wire _1400;
    wire [63:0] _1415;
    wire [63:0] _27;
    reg [63:0] _1391;
    wire [63:0] _1428;
    wire [63:0] _1424;
    wire [63:0] _1429;
    wire [63:0] _1430;
    wire _1416;
    wire [63:0] _1431;
    wire [63:0] _28;
    reg [63:0] _1411;
    wire [63:0] _1437;
    wire [63:0] _1445;
    wire [63:0] _1446;
    wire _1432;
    wire [63:0] _1447;
    wire [63:0] _29;
    reg [63:0] _1423;
    wire [63:0] _1460;
    wire [63:0] _1456;
    wire [63:0] _1461;
    wire [63:0] _1462;
    wire _1448;
    wire [63:0] _1463;
    wire [63:0] _30;
    reg [63:0] _1443;
    wire [63:0] _1469;
    wire [63:0] _1477;
    wire [63:0] _1478;
    wire _1464;
    wire [63:0] _1479;
    wire [63:0] _31;
    reg [63:0] _1455;
    wire [63:0] _1492;
    wire [63:0] _1488;
    wire [63:0] _1493;
    wire [63:0] _1494;
    wire _1480;
    wire [63:0] _1495;
    wire [63:0] _32;
    reg [63:0] _1475;
    wire [63:0] _1501;
    wire [63:0] _1509;
    wire [63:0] _1510;
    wire _1496;
    wire [63:0] _1511;
    wire [63:0] _33;
    reg [63:0] _1487;
    wire [63:0] _1524;
    wire [63:0] _1520;
    wire [63:0] _1525;
    wire [63:0] _1526;
    wire _1512;
    wire [63:0] _1527;
    wire [63:0] _34;
    reg [63:0] _1507;
    wire [63:0] _1533;
    wire [63:0] _1541;
    wire [63:0] _1542;
    wire _1528;
    wire [63:0] _1543;
    wire [63:0] _35;
    reg [63:0] _1519;
    wire [63:0] _1556;
    wire [63:0] _1552;
    wire [63:0] _1557;
    wire [63:0] _1558;
    wire _1544;
    wire [63:0] _1559;
    wire [63:0] _36;
    reg [63:0] _1539;
    wire [63:0] _1565;
    wire [63:0] _1573;
    wire [63:0] _1574;
    wire _1560;
    wire [63:0] _1575;
    wire [63:0] _37;
    reg [63:0] _1551;
    wire [63:0] _1588;
    wire [63:0] _1584;
    wire [63:0] _1589;
    wire [63:0] _1590;
    wire _1576;
    wire [63:0] _1591;
    wire [63:0] _38;
    reg [63:0] _1571;
    wire [63:0] _1597;
    wire [63:0] _1605;
    wire [63:0] _1606;
    wire _1592;
    wire [63:0] _1607;
    wire [63:0] _39;
    reg [63:0] _1583;
    wire [63:0] _1620;
    wire [63:0] _1616;
    wire [63:0] _1621;
    wire [63:0] _1622;
    wire _1608;
    wire [63:0] _1623;
    wire [63:0] _40;
    reg [63:0] _1603;
    wire [63:0] _1629;
    wire [63:0] _1637;
    wire [63:0] _1638;
    wire _1624;
    wire [63:0] _1639;
    wire [63:0] _41;
    reg [63:0] _1615;
    wire [63:0] _1652;
    wire [63:0] _1648;
    wire [63:0] _1653;
    wire [63:0] _1654;
    wire _1640;
    wire [63:0] _1655;
    wire [63:0] _42;
    reg [63:0] _1635;
    wire [63:0] _1661;
    wire [63:0] _1669;
    wire [63:0] _1670;
    wire _1656;
    wire [63:0] _1671;
    wire [63:0] _43;
    reg [63:0] _1647;
    wire [63:0] _1684;
    wire [63:0] _1680;
    wire [63:0] _1685;
    wire [63:0] _1686;
    wire _1672;
    wire [63:0] _1687;
    wire [63:0] _44;
    reg [63:0] _1667;
    wire [63:0] _1693;
    wire [63:0] _1701;
    wire [63:0] _1702;
    wire _1688;
    wire [63:0] _1703;
    wire [63:0] _45;
    reg [63:0] _1679;
    wire [63:0] _1716;
    wire [63:0] _1712;
    wire [63:0] _1717;
    wire [63:0] _1718;
    wire _1704;
    wire [63:0] _1719;
    wire [63:0] _46;
    reg [63:0] _1699;
    wire [63:0] _1725;
    wire [63:0] _1733;
    wire [63:0] _1734;
    wire _1720;
    wire [63:0] _1735;
    wire [63:0] _47;
    reg [63:0] _1711;
    wire [63:0] _1748;
    wire [63:0] _1744;
    wire [63:0] _1749;
    wire [63:0] _1750;
    wire _1736;
    wire [63:0] _1751;
    wire [63:0] _48;
    reg [63:0] _1731;
    wire [63:0] _1757;
    wire [63:0] _1765;
    wire [63:0] _1766;
    wire _1752;
    wire [63:0] _1767;
    wire [63:0] _49;
    reg [63:0] _1743;
    wire [63:0] _1780;
    wire [63:0] _1776;
    wire [63:0] _1781;
    wire [63:0] _1782;
    wire _1768;
    wire [63:0] _1783;
    wire [63:0] _50;
    reg [63:0] _1763;
    wire [63:0] _1789;
    wire [63:0] _1797;
    wire [63:0] _1798;
    wire _1784;
    wire [63:0] _1799;
    wire [63:0] _51;
    reg [63:0] _1775;
    wire [63:0] _1812;
    wire [63:0] _1808;
    wire [63:0] _1813;
    wire [63:0] _1814;
    wire _1800;
    wire [63:0] _1815;
    wire [63:0] _52;
    reg [63:0] _1795;
    wire [63:0] _1821;
    wire [63:0] _1829;
    wire [63:0] _1830;
    wire _1816;
    wire [63:0] _1831;
    wire [63:0] _53;
    reg [63:0] _1807;
    wire [63:0] _1844;
    wire [63:0] _1840;
    wire [63:0] _1845;
    wire [63:0] _1846;
    wire _1832;
    wire [63:0] _1847;
    wire [63:0] _54;
    reg [63:0] _1827;
    wire [63:0] _1853;
    wire [63:0] _1861;
    wire [63:0] _1862;
    wire _1848;
    wire [63:0] _1863;
    wire [63:0] _55;
    reg [63:0] _1839;
    wire [63:0] _1876;
    wire [63:0] _1872;
    wire [63:0] _1877;
    wire [63:0] _1878;
    wire _1864;
    wire [63:0] _1879;
    wire [63:0] _56;
    reg [63:0] _1859;
    wire [63:0] _1885;
    wire [63:0] _1893;
    wire [63:0] _1894;
    wire _1880;
    wire [63:0] _1895;
    wire [63:0] _57;
    reg [63:0] _1871;
    wire [63:0] _1908;
    wire [63:0] _1904;
    wire [63:0] _1909;
    wire [63:0] _1910;
    wire _1896;
    wire [63:0] _1911;
    wire [63:0] _58;
    reg [63:0] _1891;
    wire [63:0] _1917;
    wire [63:0] _1925;
    wire [63:0] _1926;
    wire _1912;
    wire [63:0] _1927;
    wire [63:0] _59;
    reg [63:0] _1903;
    wire [63:0] _1940;
    wire [63:0] _1936;
    wire [63:0] _1941;
    wire [63:0] _1942;
    wire _1928;
    wire [63:0] _1943;
    wire [63:0] _60;
    reg [63:0] _1923;
    wire [63:0] _1949;
    wire [63:0] _1957;
    wire [63:0] _1958;
    wire _1944;
    wire [63:0] _1959;
    wire [63:0] _61;
    reg [63:0] _1935;
    wire [63:0] _1972;
    wire [63:0] _1968;
    wire [63:0] _1973;
    wire [63:0] _1974;
    wire _1960;
    wire [63:0] _1975;
    wire [63:0] _62;
    reg [63:0] _1955;
    wire [63:0] _1981;
    wire [63:0] _1989;
    wire [63:0] _1990;
    wire _1976;
    wire [63:0] _1991;
    wire [63:0] _63;
    reg [63:0] _1967;
    wire [63:0] _2004;
    wire [63:0] _2000;
    wire [63:0] _2005;
    wire [63:0] _2006;
    wire _1992;
    wire [63:0] _2007;
    wire [63:0] _64;
    reg [63:0] _1987;
    wire [63:0] _2013;
    wire [63:0] _2021;
    wire [63:0] _2022;
    wire _2008;
    wire [63:0] _2023;
    wire [63:0] _65;
    reg [63:0] _1999;
    wire [63:0] _2036;
    wire [63:0] _2032;
    wire [63:0] _2037;
    wire [63:0] _2038;
    wire _2024;
    wire [63:0] _2039;
    wire [63:0] _66;
    reg [63:0] _2019;
    wire [63:0] _2045;
    wire [63:0] _2053;
    wire [63:0] _2054;
    wire _2040;
    wire [63:0] _2055;
    wire [63:0] _67;
    reg [63:0] _2031;
    wire [63:0] _2068;
    wire [63:0] _2064;
    wire [63:0] _2069;
    wire [63:0] _2070;
    wire _2056;
    wire [63:0] _2071;
    wire [63:0] _68;
    reg [63:0] _2051;
    wire [63:0] _2077;
    wire [63:0] _2085;
    wire [63:0] _2086;
    wire _2072;
    wire [63:0] _2087;
    wire [63:0] _69;
    reg [63:0] _2063;
    wire [63:0] _2100;
    wire [63:0] _2096;
    wire [63:0] _2101;
    wire [63:0] _2102;
    wire _2088;
    wire [63:0] _2103;
    wire [63:0] _70;
    reg [63:0] _2083;
    wire [63:0] _2109;
    wire [63:0] _2117;
    wire [63:0] _2118;
    wire _2104;
    wire [63:0] _2119;
    wire [63:0] _71;
    reg [63:0] _2095;
    wire [63:0] _2132;
    wire [63:0] _2128;
    wire [63:0] _2133;
    wire [63:0] _2134;
    wire _2120;
    wire [63:0] _2135;
    wire [63:0] _72;
    reg [63:0] _2115;
    wire [63:0] _2141;
    wire [63:0] _2149;
    wire [63:0] _2150;
    wire _2136;
    wire [63:0] _2151;
    wire [63:0] _73;
    reg [63:0] _2127;
    wire [63:0] _2164;
    wire [63:0] _2160;
    wire [63:0] _2165;
    wire [63:0] _2166;
    wire _2152;
    wire [63:0] _2167;
    wire [63:0] _74;
    reg [63:0] _2147;
    wire [63:0] _2173;
    wire [63:0] _2181;
    wire [63:0] _2182;
    wire _2168;
    wire [63:0] _2183;
    wire [63:0] _75;
    reg [63:0] _2159;
    wire [63:0] _2196;
    wire [63:0] _2192;
    wire [63:0] _2197;
    wire [63:0] _2198;
    wire _2184;
    wire [63:0] _2199;
    wire [63:0] _76;
    reg [63:0] _2179;
    wire [63:0] _2205;
    wire [63:0] _2213;
    wire [63:0] _2214;
    wire _2200;
    wire [63:0] _2215;
    wire [63:0] _77;
    reg [63:0] _2191;
    wire [63:0] _2228;
    wire [63:0] _2224;
    wire [63:0] _2229;
    wire [63:0] _2230;
    wire _2216;
    wire [63:0] _2231;
    wire [63:0] _78;
    reg [63:0] _2211;
    wire [63:0] _2237;
    wire [63:0] _2245;
    wire [63:0] _2246;
    wire _2232;
    wire [63:0] _2247;
    wire [63:0] _79;
    reg [63:0] _2223;
    wire [63:0] _2260;
    wire [63:0] _2256;
    wire [63:0] _2261;
    wire [63:0] _2262;
    wire _2248;
    wire [63:0] _2263;
    wire [63:0] _80;
    reg [63:0] _2243;
    wire [63:0] _2269;
    wire [63:0] _2277;
    wire [63:0] _2278;
    wire _2264;
    wire [63:0] _2279;
    wire [63:0] _81;
    reg [63:0] _2255;
    wire [63:0] _2292;
    wire [63:0] _2288;
    wire [63:0] _2293;
    wire [63:0] _2294;
    wire _2280;
    wire [63:0] _2295;
    wire [63:0] _82;
    reg [63:0] _2275;
    wire [63:0] _2301;
    wire [63:0] _2309;
    wire [63:0] _2310;
    wire _2296;
    wire [63:0] _2311;
    wire [63:0] _83;
    reg [63:0] _2287;
    wire [63:0] _2324;
    wire [63:0] _2320;
    wire [63:0] _2325;
    wire [63:0] _2326;
    wire _2312;
    wire [63:0] _2327;
    wire [63:0] _84;
    reg [63:0] _2307;
    wire [63:0] _2333;
    wire [63:0] _2341;
    wire [63:0] _2342;
    wire _2328;
    wire [63:0] _2343;
    wire [63:0] _85;
    reg [63:0] _2319;
    wire [63:0] _2356;
    wire [63:0] _2352;
    wire [63:0] _2357;
    wire [63:0] _2358;
    wire _2344;
    wire [63:0] _2359;
    wire [63:0] _86;
    reg [63:0] _2339;
    wire [63:0] _2365;
    wire [63:0] _2373;
    wire [63:0] _2374;
    wire _2360;
    wire [63:0] _2375;
    wire [63:0] _87;
    reg [63:0] _2351;
    wire [63:0] _2388;
    wire [63:0] _2384;
    wire [63:0] _2389;
    wire [63:0] _2390;
    wire _2376;
    wire [63:0] _2391;
    wire [63:0] _88;
    reg [63:0] _2371;
    wire [63:0] _2397;
    wire [63:0] _2405;
    wire [63:0] _2406;
    wire _2392;
    wire [63:0] _2407;
    wire [63:0] _89;
    reg [63:0] _2383;
    wire [63:0] _2420;
    wire [63:0] _2416;
    wire [63:0] _2421;
    wire [63:0] _2422;
    wire _2408;
    wire [63:0] _2423;
    wire [63:0] _90;
    reg [63:0] _2403;
    wire [63:0] _2429;
    wire [63:0] _2437;
    wire [63:0] _2438;
    wire _2424;
    wire [63:0] _2439;
    wire [63:0] _91;
    reg [63:0] _2415;
    wire [63:0] _2452;
    wire [63:0] _2448;
    wire [63:0] _2453;
    wire [63:0] _2454;
    wire _2440;
    wire [63:0] _2455;
    wire [63:0] _92;
    reg [63:0] _2435;
    wire [63:0] _2461;
    wire [63:0] _2469;
    wire [63:0] _2470;
    wire _2456;
    wire [63:0] _2471;
    wire [63:0] _93;
    reg [63:0] _2447;
    wire [63:0] _2484;
    wire [63:0] _2480;
    wire [63:0] _2485;
    wire [63:0] _2486;
    wire _2472;
    wire [63:0] _2487;
    wire [63:0] _94;
    reg [63:0] _2467;
    wire [63:0] _2493;
    wire [63:0] _2501;
    wire [63:0] _2502;
    wire _2488;
    wire [63:0] _2503;
    wire [63:0] _95;
    reg [63:0] _2479;
    wire [63:0] _2516;
    wire [63:0] _2512;
    wire [63:0] _2517;
    wire [63:0] _2518;
    wire _2504;
    wire [63:0] _2519;
    wire [63:0] _96;
    reg [63:0] _2499;
    wire [63:0] _2525;
    wire [63:0] _2533;
    wire [63:0] _2534;
    wire _2520;
    wire [63:0] _2535;
    wire [63:0] _97;
    reg [63:0] _2511;
    wire [63:0] _2548;
    wire [63:0] _2544;
    wire [63:0] _2549;
    wire [63:0] _2550;
    wire _2536;
    wire [63:0] _2551;
    wire [63:0] _98;
    reg [63:0] _2531;
    wire [63:0] _2557;
    wire [63:0] _2565;
    wire [63:0] _2566;
    wire _2552;
    wire [63:0] _2567;
    wire [63:0] _99;
    reg [63:0] _2543;
    wire [63:0] _2580;
    wire [63:0] _2576;
    wire [63:0] _2581;
    wire [63:0] _2582;
    wire _2568;
    wire [63:0] _2583;
    wire [63:0] _100;
    reg [63:0] _2563;
    wire [63:0] _2589;
    wire [63:0] _2597;
    wire [63:0] _2598;
    wire _2584;
    wire [63:0] _2599;
    wire [63:0] _101;
    reg [63:0] _2575;
    wire [63:0] _2612;
    wire [63:0] _2608;
    wire [63:0] _2613;
    wire [63:0] _2614;
    wire _2600;
    wire [63:0] _2615;
    wire [63:0] _102;
    reg [63:0] _2595;
    wire [63:0] _2621;
    wire [63:0] _2629;
    wire [63:0] _2630;
    wire _2616;
    wire [63:0] _2631;
    wire [63:0] _103;
    reg [63:0] _2607;
    wire [63:0] _2644;
    wire [63:0] _2640;
    wire [63:0] _2645;
    wire [63:0] _2646;
    wire _2632;
    wire [63:0] _2647;
    wire [63:0] _104;
    reg [63:0] _2627;
    wire [63:0] _2653;
    wire [63:0] _2661;
    wire [63:0] _2662;
    wire _2648;
    wire [63:0] _2663;
    wire [63:0] _105;
    reg [63:0] _2639;
    wire [63:0] _2676;
    wire [63:0] _2672;
    wire [63:0] _2677;
    wire [63:0] _2678;
    wire _2664;
    wire [63:0] _2679;
    wire [63:0] _106;
    reg [63:0] _2659;
    wire [63:0] _2685;
    wire [63:0] _2693;
    wire [63:0] _2694;
    wire _2680;
    wire [63:0] _2695;
    wire [63:0] _107;
    reg [63:0] _2671;
    wire [63:0] _2708;
    wire [63:0] _2704;
    wire [63:0] _2709;
    wire [63:0] _2710;
    wire _2696;
    wire [63:0] _2711;
    wire [63:0] _108;
    reg [63:0] _2691;
    wire [63:0] _2717;
    wire [63:0] _2725;
    wire [63:0] _2726;
    wire _2712;
    wire [63:0] _2727;
    wire [63:0] _109;
    reg [63:0] _2703;
    wire [63:0] _2740;
    wire [63:0] _2736;
    wire [63:0] _2741;
    wire [63:0] _2742;
    wire _2728;
    wire [63:0] _2743;
    wire [63:0] _110;
    reg [63:0] _2723;
    wire [63:0] _2749;
    wire [63:0] _2757;
    wire [63:0] _2758;
    wire _2744;
    wire [63:0] _2759;
    wire [63:0] _111;
    reg [63:0] _2735;
    wire [63:0] _2772;
    wire [63:0] _2768;
    wire [63:0] _2773;
    wire [63:0] _2774;
    wire _2760;
    wire [63:0] _2775;
    wire [63:0] _112;
    reg [63:0] _2755;
    wire [63:0] _2781;
    wire [63:0] _2789;
    wire [63:0] _2790;
    wire _2776;
    wire [63:0] _2791;
    wire [63:0] _113;
    reg [63:0] _2767;
    wire [63:0] _2804;
    wire [63:0] _2800;
    wire [63:0] _2805;
    wire [63:0] _2806;
    wire _2792;
    wire [63:0] _2807;
    wire [63:0] _114;
    reg [63:0] _2787;
    wire [63:0] _2813;
    wire [63:0] _2821;
    wire [63:0] _2822;
    wire _2808;
    wire [63:0] _2823;
    wire [63:0] _115;
    reg [63:0] _2799;
    wire [63:0] _2836;
    wire [63:0] _2832;
    wire [63:0] _2837;
    wire [63:0] _2838;
    wire _2824;
    wire [63:0] _2839;
    wire [63:0] _116;
    reg [63:0] _2819;
    wire [63:0] _2845;
    wire [63:0] _2853;
    wire [63:0] _2854;
    wire _2840;
    wire [63:0] _2855;
    wire [63:0] _117;
    reg [63:0] _2831;
    wire [63:0] _2868;
    wire [63:0] _2864;
    wire [63:0] _2869;
    wire [63:0] _2870;
    wire _2856;
    wire [63:0] _2871;
    wire [63:0] _118;
    reg [63:0] _2851;
    wire [63:0] _2877;
    wire [63:0] _2885;
    wire [63:0] _2886;
    wire _2872;
    wire [63:0] _2887;
    wire [63:0] _119;
    reg [63:0] _2863;
    wire [63:0] _2900;
    wire [63:0] _2896;
    wire [63:0] _2901;
    wire [63:0] _2902;
    wire _2888;
    wire [63:0] _2903;
    wire [63:0] _120;
    reg [63:0] _2883;
    wire [63:0] _2909;
    wire [63:0] _2917;
    wire [63:0] _2918;
    wire _2904;
    wire [63:0] _2919;
    wire [63:0] _121;
    reg [63:0] _2895;
    wire [63:0] _2932;
    wire [63:0] _2928;
    wire [63:0] _2933;
    wire [63:0] _2934;
    wire _2920;
    wire [63:0] _2935;
    wire [63:0] _122;
    reg [63:0] _2915;
    wire [63:0] _2941;
    wire [63:0] _2949;
    wire [63:0] _2950;
    wire _2936;
    wire [63:0] _2951;
    wire [63:0] _123;
    reg [63:0] _2927;
    wire [63:0] _2964;
    wire [63:0] _2960;
    wire [63:0] _2965;
    wire [63:0] _2966;
    wire _2952;
    wire [63:0] _2967;
    wire [63:0] _124;
    reg [63:0] _2947;
    wire [63:0] _2973;
    wire [63:0] _2981;
    wire [63:0] _2982;
    wire _2968;
    wire [63:0] _2983;
    wire [63:0] _125;
    reg [63:0] _2959;
    wire [63:0] _2996;
    wire [63:0] _2992;
    wire [63:0] _2997;
    wire [63:0] _2998;
    wire _2984;
    wire [63:0] _2999;
    wire [63:0] _126;
    reg [63:0] _2979;
    wire [63:0] _3005;
    wire [63:0] _3013;
    wire [63:0] _3014;
    wire _3000;
    wire [63:0] _3015;
    wire [63:0] _127;
    reg [63:0] _2991;
    wire [63:0] _3028;
    wire [63:0] _3024;
    wire [63:0] _3029;
    wire [63:0] _3030;
    wire _3016;
    wire [63:0] _3031;
    wire [63:0] _128;
    reg [63:0] _3011;
    wire [63:0] _3037;
    wire [63:0] _3045;
    wire [63:0] _3046;
    wire _3032;
    wire [63:0] _3047;
    wire [63:0] _129;
    reg [63:0] _3023;
    wire [63:0] _3060;
    wire [63:0] _3056;
    wire [63:0] _3061;
    wire [63:0] _3062;
    wire _3048;
    wire [63:0] _3063;
    wire [63:0] _130;
    reg [63:0] _3043;
    wire [63:0] _3069;
    wire [63:0] _3077;
    wire [63:0] _3078;
    wire _3064;
    wire [63:0] _3079;
    wire [63:0] _131;
    reg [63:0] _3055;
    wire [63:0] _3092;
    wire [63:0] _3088;
    wire [63:0] _3093;
    wire [63:0] _3094;
    wire _3080;
    wire [63:0] _3095;
    wire [63:0] _132;
    reg [63:0] _3075;
    wire [63:0] _3101;
    wire [63:0] _3109;
    wire [63:0] _3110;
    wire _3096;
    wire [63:0] _3111;
    wire [63:0] _133;
    reg [63:0] _3087;
    wire [63:0] _3124;
    wire [63:0] _3120;
    wire [63:0] _3125;
    wire [63:0] _3126;
    wire _3112;
    wire [63:0] _3127;
    wire [63:0] _134;
    reg [63:0] _3107;
    wire [63:0] _3133;
    wire [63:0] _3141;
    wire [63:0] _3142;
    wire _3128;
    wire [63:0] _3143;
    wire [63:0] _135;
    reg [63:0] _3119;
    wire [63:0] _3156;
    wire [63:0] _3152;
    wire [63:0] _3157;
    wire [63:0] _3158;
    wire _3144;
    wire [63:0] _3159;
    wire [63:0] _136;
    reg [63:0] _3139;
    wire [63:0] _3165;
    wire [63:0] _3173;
    wire [63:0] _3174;
    wire _3160;
    wire [63:0] _3175;
    wire [63:0] _137;
    reg [63:0] _3151;
    wire [63:0] _3188;
    wire [63:0] _3184;
    wire [63:0] _3189;
    wire [63:0] _3190;
    wire _3176;
    wire [63:0] _3191;
    wire [63:0] _138;
    reg [63:0] _3171;
    wire [63:0] _3197;
    wire [63:0] _3205;
    wire [63:0] _3206;
    wire _3192;
    wire [63:0] _3207;
    wire [63:0] _139;
    reg [63:0] _3183;
    wire [63:0] _3220;
    wire [63:0] _3216;
    wire [63:0] _3221;
    wire [63:0] _3222;
    wire _3208;
    wire [63:0] _3223;
    wire [63:0] _140;
    reg [63:0] _3203;
    wire [63:0] _3229;
    wire [63:0] _3237;
    wire [63:0] _3238;
    wire _3224;
    wire [63:0] _3239;
    wire [63:0] _141;
    reg [63:0] _3215;
    wire [63:0] _3252;
    wire [63:0] _3248;
    wire [63:0] _3253;
    wire [63:0] _3254;
    wire _3240;
    wire [63:0] _3255;
    wire [63:0] _142;
    reg [63:0] _3235;
    wire [63:0] _3261;
    wire [63:0] _3269;
    wire [63:0] _3270;
    wire _3256;
    wire [63:0] _3271;
    wire [63:0] _143;
    reg [63:0] _3247;
    wire [63:0] _3284;
    wire [63:0] _3280;
    wire [63:0] _3285;
    wire [63:0] _3286;
    wire _3272;
    wire [63:0] _3287;
    wire [63:0] _144;
    reg [63:0] _3267;
    wire [63:0] _3293;
    wire [63:0] _3301;
    wire [63:0] _3302;
    wire _3288;
    wire [63:0] _3303;
    wire [63:0] _145;
    reg [63:0] _3279;
    wire [63:0] _3316;
    wire [63:0] _3312;
    wire [63:0] _3317;
    wire [63:0] _3318;
    wire _3304;
    wire [63:0] _3319;
    wire [63:0] _146;
    reg [63:0] _3299;
    wire [63:0] _3325;
    wire [63:0] _3333;
    wire [63:0] _3334;
    wire _3320;
    wire [63:0] _3335;
    wire [63:0] _147;
    reg [63:0] _3311;
    wire [63:0] _3348;
    wire [63:0] _3344;
    wire [63:0] _3349;
    wire [63:0] _3350;
    wire _3336;
    wire [63:0] _3351;
    wire [63:0] _148;
    reg [63:0] _3331;
    wire [63:0] _3357;
    wire [63:0] _3365;
    wire [63:0] _3366;
    wire _3352;
    wire [63:0] _3367;
    wire [63:0] _149;
    reg [63:0] _3343;
    wire [63:0] _3380;
    wire [63:0] _3376;
    wire [63:0] _3381;
    wire [63:0] _3382;
    wire _3368;
    wire [63:0] _3383;
    wire [63:0] _150;
    reg [63:0] _3363;
    wire [63:0] _3389;
    wire [63:0] _3397;
    wire [63:0] _3398;
    wire _3384;
    wire [63:0] _3399;
    wire [63:0] _151;
    reg [63:0] _3375;
    wire [63:0] _3412;
    wire [63:0] _3408;
    wire [63:0] _3413;
    wire [63:0] _3414;
    wire _3400;
    wire [63:0] _3415;
    wire [63:0] _152;
    reg [63:0] _3395;
    wire [63:0] _3421;
    wire [63:0] _3429;
    wire [63:0] _3430;
    wire _3416;
    wire [63:0] _3431;
    wire [63:0] _153;
    reg [63:0] _3407;
    wire [63:0] _3444;
    wire [63:0] _3440;
    wire [63:0] _3445;
    wire [63:0] _3446;
    wire _3432;
    wire [63:0] _3447;
    wire [63:0] _154;
    reg [63:0] _3427;
    wire [63:0] _3453;
    wire [63:0] _3461;
    wire [63:0] _3462;
    wire _3448;
    wire [63:0] _3463;
    wire [63:0] _155;
    reg [63:0] _3439;
    wire [63:0] _3476;
    wire [63:0] _3472;
    wire [63:0] _3477;
    wire [63:0] _3478;
    wire _3464;
    wire [63:0] _3479;
    wire [63:0] _156;
    reg [63:0] _3459;
    wire [63:0] _3485;
    wire [63:0] _3493;
    wire [63:0] _3494;
    wire _3480;
    wire [63:0] _3495;
    wire [63:0] _157;
    reg [63:0] _3471;
    wire [63:0] _3508;
    wire [63:0] _3504;
    wire [63:0] _3509;
    wire [63:0] _3510;
    wire _3496;
    wire [63:0] _3511;
    wire [63:0] _158;
    reg [63:0] _3491;
    wire [63:0] _3517;
    wire [63:0] _3525;
    wire [63:0] _3526;
    wire _3512;
    wire [63:0] _3527;
    wire [63:0] _159;
    reg [63:0] _3503;
    wire [63:0] _3540;
    wire [63:0] _3536;
    wire [63:0] _3541;
    wire [63:0] _3542;
    wire _3528;
    wire [63:0] _3543;
    wire [63:0] _160;
    reg [63:0] _3523;
    wire [63:0] _3549;
    wire [63:0] _3557;
    wire [63:0] _3558;
    wire _3544;
    wire [63:0] _3559;
    wire [63:0] _161;
    reg [63:0] _3535;
    wire [63:0] _3572;
    wire [63:0] _3568;
    wire [63:0] _3573;
    wire [63:0] _3574;
    wire _3560;
    wire [63:0] _3575;
    wire [63:0] _162;
    reg [63:0] _3555;
    wire [63:0] _3581;
    wire [63:0] _3589;
    wire [63:0] _3590;
    wire _3576;
    wire [63:0] _3591;
    wire [63:0] _163;
    reg [63:0] _3567;
    wire [63:0] _3604;
    wire [63:0] _3600;
    wire [63:0] _3605;
    wire [63:0] _3606;
    wire _3592;
    wire [63:0] _3607;
    wire [63:0] _164;
    reg [63:0] _3587;
    wire [63:0] _3613;
    wire [63:0] _3621;
    wire [63:0] _3622;
    wire _3608;
    wire [63:0] _3623;
    wire [63:0] _165;
    reg [63:0] _3599;
    wire [63:0] _3636;
    wire [63:0] _3632;
    wire [63:0] _3637;
    wire [63:0] _3638;
    wire _3624;
    wire [63:0] _3639;
    wire [63:0] _166;
    reg [63:0] _3619;
    wire [63:0] _3645;
    wire [63:0] _3653;
    wire [63:0] _3654;
    wire _3640;
    wire [63:0] _3655;
    wire [63:0] _167;
    reg [63:0] _3631;
    wire [63:0] _3668;
    wire [63:0] _3664;
    wire [63:0] _3669;
    wire [63:0] _3670;
    wire _3656;
    wire [63:0] _3671;
    wire [63:0] _168;
    reg [63:0] _3651;
    wire [63:0] _3677;
    wire [63:0] _3685;
    wire [63:0] _3686;
    wire _3672;
    wire [63:0] _3687;
    wire [63:0] _169;
    reg [63:0] _3663;
    wire [63:0] _3700;
    wire [63:0] _3696;
    wire [63:0] _3701;
    wire [63:0] _3702;
    wire _3688;
    wire [63:0] _3703;
    wire [63:0] _170;
    reg [63:0] _3683;
    wire [63:0] _3709;
    wire [63:0] _3717;
    wire [63:0] _3718;
    wire _3704;
    wire [63:0] _3719;
    wire [63:0] _171;
    reg [63:0] _3695;
    wire [63:0] _3732;
    wire [63:0] _3728;
    wire [63:0] _3733;
    wire [63:0] _3734;
    wire _3720;
    wire [63:0] _3735;
    wire [63:0] _172;
    reg [63:0] _3715;
    wire [63:0] _3741;
    wire [63:0] _3749;
    wire [63:0] _3750;
    wire _3736;
    wire [63:0] _3751;
    wire [63:0] _173;
    reg [63:0] _3727;
    wire [63:0] _3764;
    wire [63:0] _3760;
    wire [63:0] _3765;
    wire [63:0] _3766;
    wire _3752;
    wire [63:0] _3767;
    wire [63:0] _174;
    reg [63:0] _3747;
    wire [63:0] _3773;
    wire [63:0] _3781;
    wire [63:0] _3782;
    wire _3768;
    wire [63:0] _3783;
    wire [63:0] _175;
    reg [63:0] _3759;
    wire [63:0] _3796;
    wire [63:0] _3792;
    wire [63:0] _3797;
    wire [63:0] _3798;
    wire _3784;
    wire [63:0] _3799;
    wire [63:0] _176;
    reg [63:0] _3779;
    wire [63:0] _3805;
    wire [63:0] _3813;
    wire [63:0] _3814;
    wire _3800;
    wire [63:0] _3815;
    wire [63:0] _177;
    reg [63:0] _3791;
    wire [63:0] _3828;
    wire [63:0] _3824;
    wire [63:0] _3829;
    wire [63:0] _3830;
    wire _3816;
    wire [63:0] _3831;
    wire [63:0] _178;
    reg [63:0] _3811;
    wire [63:0] _3837;
    wire [63:0] _3845;
    wire [63:0] _3846;
    wire _3832;
    wire [63:0] _3847;
    wire [63:0] _179;
    reg [63:0] _3823;
    wire [63:0] _3860;
    wire [63:0] _3856;
    wire [63:0] _3861;
    wire [63:0] _3862;
    wire _3848;
    wire [63:0] _3863;
    wire [63:0] _180;
    reg [63:0] _3843;
    wire [63:0] _3869;
    wire [63:0] _3877;
    wire [63:0] _3878;
    wire _3864;
    wire [63:0] _3879;
    wire [63:0] _181;
    reg [63:0] _3855;
    wire [63:0] _3892;
    wire [63:0] _3888;
    wire [63:0] _3893;
    wire [63:0] _3894;
    wire _3880;
    wire [63:0] _3895;
    wire [63:0] _182;
    reg [63:0] _3875;
    wire [63:0] _3901;
    wire [63:0] _3909;
    wire [63:0] _3910;
    wire _3896;
    wire [63:0] _3911;
    wire [63:0] _183;
    reg [63:0] _3887;
    wire [63:0] _3924;
    wire [63:0] _3920;
    wire [63:0] _3925;
    wire [63:0] _3926;
    wire _3912;
    wire [63:0] _3927;
    wire [63:0] _184;
    reg [63:0] _3907;
    wire [63:0] _3933;
    wire [63:0] _3941;
    wire [63:0] _3942;
    wire _3928;
    wire [63:0] _3943;
    wire [63:0] _185;
    reg [63:0] _3919;
    wire [63:0] _3956;
    wire [63:0] _3952;
    wire [63:0] _3957;
    wire [63:0] _3958;
    wire _3944;
    wire [63:0] _3959;
    wire [63:0] _186;
    reg [63:0] _3939;
    wire [63:0] _3965;
    wire [63:0] _3973;
    wire [63:0] _3974;
    wire _3960;
    wire [63:0] _3975;
    wire [63:0] _187;
    reg [63:0] _3951;
    wire [63:0] _3988;
    wire [63:0] _3984;
    wire [63:0] _3989;
    wire [63:0] _3990;
    wire _3976;
    wire [63:0] _3991;
    wire [63:0] _188;
    reg [63:0] _3971;
    wire [63:0] _3997;
    wire [63:0] _4005;
    wire [63:0] _4006;
    wire _3992;
    wire [63:0] _4007;
    wire [63:0] _189;
    reg [63:0] _3983;
    wire [63:0] _4020;
    wire [63:0] _4016;
    wire [63:0] _4021;
    wire [63:0] _4022;
    wire _4008;
    wire [63:0] _4023;
    wire [63:0] _190;
    reg [63:0] _4003;
    wire [63:0] _4029;
    wire [63:0] _4037;
    wire [63:0] _4038;
    wire _4024;
    wire [63:0] _4039;
    wire [63:0] _191;
    reg [63:0] _4015;
    wire [63:0] _4052;
    wire [63:0] _4048;
    wire [63:0] _4053;
    wire [63:0] _4054;
    wire _4040;
    wire [63:0] _4055;
    wire [63:0] _192;
    reg [63:0] _4035;
    wire [63:0] _4061;
    wire [63:0] _4069;
    wire [63:0] _4070;
    wire _4056;
    wire [63:0] _4071;
    wire [63:0] _193;
    reg [63:0] _4047;
    wire [63:0] _4084;
    wire [63:0] _4080;
    wire [63:0] _4085;
    wire [63:0] _4086;
    wire _4072;
    wire [63:0] _4087;
    wire [63:0] _194;
    reg [63:0] _4067;
    wire [63:0] _4093;
    wire [63:0] _4101;
    wire [63:0] _4102;
    wire _4088;
    wire [63:0] _4103;
    wire [63:0] _195;
    reg [63:0] _4079;
    wire [63:0] _4116;
    wire [63:0] _4112;
    wire [63:0] _4117;
    wire [63:0] _4118;
    wire _4104;
    wire [63:0] _4119;
    wire [63:0] _196;
    reg [63:0] _4099;
    wire [63:0] _4125;
    wire [63:0] _4133;
    wire [63:0] _4134;
    wire _4120;
    wire [63:0] _4135;
    wire [63:0] _197;
    reg [63:0] _4111;
    wire [63:0] _4148;
    wire [63:0] _4144;
    wire [63:0] _4149;
    wire [63:0] _4150;
    wire _4136;
    wire [63:0] _4151;
    wire [63:0] _198;
    reg [63:0] _4131;
    wire [63:0] _4157;
    wire [63:0] _4165;
    wire [63:0] _4166;
    wire _4152;
    wire [63:0] _4167;
    wire [63:0] _199;
    reg [63:0] _4143;
    wire [63:0] _4180;
    wire [63:0] _4176;
    wire [63:0] _4181;
    wire [63:0] _4182;
    wire _4168;
    wire [63:0] _4183;
    wire [63:0] _200;
    reg [63:0] _4163;
    wire [63:0] _4189;
    wire [63:0] _4197;
    wire [63:0] _4198;
    wire _4184;
    wire [63:0] _4199;
    wire [63:0] _201;
    reg [63:0] _4175;
    wire [63:0] _4212;
    wire [63:0] _4208;
    wire [63:0] _4213;
    wire [63:0] _4214;
    wire _4200;
    wire [63:0] _4215;
    wire [63:0] _202;
    reg [63:0] _4195;
    wire [63:0] _4221;
    wire [63:0] _4229;
    wire [63:0] _4230;
    wire _4216;
    wire [63:0] _4231;
    wire [63:0] _203;
    reg [63:0] _4207;
    wire [63:0] _4244;
    wire [63:0] _4240;
    wire [63:0] _4245;
    wire [63:0] _4246;
    wire _4232;
    wire [63:0] _4247;
    wire [63:0] _204;
    reg [63:0] _4227;
    wire [64:0] _5439;
    wire [64:0] _4242;
    wire [64:0] _4223;
    wire [64:0] _4222;
    wire _4224;
    wire [63:0] _5432;
    wire [64:0] _4219;
    wire [64:0] _4210;
    wire [64:0] _4191;
    wire [64:0] _4190;
    wire _4192;
    wire [63:0] _5420;
    wire [64:0] _4187;
    wire [64:0] _4178;
    wire [64:0] _4159;
    wire [64:0] _4158;
    wire _4160;
    wire [63:0] _5408;
    wire [64:0] _4155;
    wire [64:0] _4146;
    wire [64:0] _4127;
    wire [64:0] _4126;
    wire _4128;
    wire [63:0] _5396;
    wire [64:0] _4123;
    wire [64:0] _4114;
    wire [64:0] _4095;
    wire [64:0] _4094;
    wire _4096;
    wire [63:0] _5384;
    wire [64:0] _4091;
    wire [64:0] _4082;
    wire [64:0] _4063;
    wire [64:0] _4062;
    wire _4064;
    wire [63:0] _5372;
    wire [64:0] _4059;
    wire [64:0] _4050;
    wire [64:0] _4031;
    wire [64:0] _4030;
    wire _4032;
    wire [63:0] _5360;
    wire [64:0] _4027;
    wire [64:0] _4018;
    wire [64:0] _3999;
    wire [64:0] _3998;
    wire _4000;
    wire [63:0] _5348;
    wire [64:0] _3995;
    wire [64:0] _3986;
    wire [64:0] _3967;
    wire [64:0] _3966;
    wire _3968;
    wire [63:0] _5336;
    wire [64:0] _3963;
    wire [64:0] _3954;
    wire [64:0] _3935;
    wire [64:0] _3934;
    wire _3936;
    wire [63:0] _5324;
    wire [64:0] _3931;
    wire [64:0] _3922;
    wire [64:0] _3903;
    wire [64:0] _3902;
    wire _3904;
    wire [63:0] _5312;
    wire [64:0] _3899;
    wire [64:0] _3890;
    wire [64:0] _3871;
    wire [64:0] _3870;
    wire _3872;
    wire [63:0] _5300;
    wire [64:0] _3867;
    wire [64:0] _3858;
    wire [64:0] _3839;
    wire [64:0] _3838;
    wire _3840;
    wire [63:0] _5288;
    wire [64:0] _3835;
    wire [64:0] _3826;
    wire [64:0] _3807;
    wire [64:0] _3806;
    wire _3808;
    wire [63:0] _5276;
    wire [64:0] _3803;
    wire [64:0] _3794;
    wire [64:0] _3775;
    wire [64:0] _3774;
    wire _3776;
    wire [63:0] _5264;
    wire [64:0] _3771;
    wire [64:0] _3762;
    wire [64:0] _3743;
    wire [64:0] _3742;
    wire _3744;
    wire [63:0] _5252;
    wire [64:0] _3739;
    wire [64:0] _3730;
    wire [64:0] _3711;
    wire [64:0] _3710;
    wire _3712;
    wire [63:0] _5240;
    wire [64:0] _3707;
    wire [64:0] _3698;
    wire [64:0] _3679;
    wire [64:0] _3678;
    wire _3680;
    wire [63:0] _5228;
    wire [64:0] _3675;
    wire [64:0] _3666;
    wire [64:0] _3647;
    wire [64:0] _3646;
    wire _3648;
    wire [63:0] _5216;
    wire [64:0] _3643;
    wire [64:0] _3634;
    wire [64:0] _3615;
    wire [64:0] _3614;
    wire _3616;
    wire [63:0] _5204;
    wire [64:0] _3611;
    wire [64:0] _3602;
    wire [64:0] _3583;
    wire [64:0] _3582;
    wire _3584;
    wire [63:0] _5192;
    wire [64:0] _3579;
    wire [64:0] _3570;
    wire [64:0] _3551;
    wire [64:0] _3550;
    wire _3552;
    wire [63:0] _5180;
    wire [64:0] _3547;
    wire [64:0] _3538;
    wire [64:0] _3519;
    wire [64:0] _3518;
    wire _3520;
    wire [63:0] _5168;
    wire [64:0] _3515;
    wire [64:0] _3506;
    wire [64:0] _3487;
    wire [64:0] _3486;
    wire _3488;
    wire [63:0] _5156;
    wire [64:0] _3483;
    wire [64:0] _3474;
    wire [64:0] _3455;
    wire [64:0] _3454;
    wire _3456;
    wire [63:0] _5144;
    wire [64:0] _3451;
    wire [64:0] _3442;
    wire [64:0] _3423;
    wire [64:0] _3422;
    wire _3424;
    wire [63:0] _5132;
    wire [64:0] _3419;
    wire [64:0] _3410;
    wire [64:0] _3391;
    wire [64:0] _3390;
    wire _3392;
    wire [63:0] _5120;
    wire [64:0] _3387;
    wire [64:0] _3378;
    wire [64:0] _3359;
    wire [64:0] _3358;
    wire _3360;
    wire [63:0] _5108;
    wire [64:0] _3355;
    wire [64:0] _3346;
    wire [64:0] _3327;
    wire [64:0] _3326;
    wire _3328;
    wire [63:0] _5096;
    wire [64:0] _3323;
    wire [64:0] _3314;
    wire [64:0] _3295;
    wire [64:0] _3294;
    wire _3296;
    wire [63:0] _5084;
    wire [64:0] _3291;
    wire [64:0] _3282;
    wire [64:0] _3263;
    wire [64:0] _3262;
    wire _3264;
    wire [63:0] _5072;
    wire [64:0] _3259;
    wire [64:0] _3250;
    wire [64:0] _3231;
    wire [64:0] _3230;
    wire _3232;
    wire [63:0] _5060;
    wire [64:0] _3227;
    wire [64:0] _3218;
    wire [64:0] _3199;
    wire [64:0] _3198;
    wire _3200;
    wire [63:0] _5048;
    wire [64:0] _3195;
    wire [64:0] _3186;
    wire [64:0] _3167;
    wire [64:0] _3166;
    wire _3168;
    wire [63:0] _5036;
    wire [64:0] _3163;
    wire [64:0] _3154;
    wire [64:0] _3135;
    wire [64:0] _3134;
    wire _3136;
    wire [63:0] _5024;
    wire [64:0] _3131;
    wire [64:0] _3122;
    wire [64:0] _3103;
    wire [64:0] _3102;
    wire _3104;
    wire [63:0] _5012;
    wire [64:0] _3099;
    wire [64:0] _3090;
    wire [64:0] _3071;
    wire [64:0] _3070;
    wire _3072;
    wire [63:0] _5000;
    wire [64:0] _3067;
    wire [64:0] _3058;
    wire [64:0] _3039;
    wire [64:0] _3038;
    wire _3040;
    wire [63:0] _4988;
    wire [64:0] _3035;
    wire [64:0] _3026;
    wire [64:0] _3007;
    wire [64:0] _3006;
    wire _3008;
    wire [63:0] _4976;
    wire [64:0] _3003;
    wire [64:0] _2994;
    wire [64:0] _2975;
    wire [64:0] _2974;
    wire _2976;
    wire [63:0] _4964;
    wire [64:0] _2971;
    wire [64:0] _2962;
    wire [64:0] _2943;
    wire [64:0] _2942;
    wire _2944;
    wire [63:0] _4952;
    wire [64:0] _2939;
    wire [64:0] _2930;
    wire [64:0] _2911;
    wire [64:0] _2910;
    wire _2912;
    wire [63:0] _4940;
    wire [64:0] _2907;
    wire [64:0] _2898;
    wire [64:0] _2879;
    wire [64:0] _2878;
    wire _2880;
    wire [63:0] _4928;
    wire [64:0] _2875;
    wire [64:0] _2866;
    wire [64:0] _2847;
    wire [64:0] _2846;
    wire _2848;
    wire [63:0] _4916;
    wire [64:0] _2843;
    wire [64:0] _2834;
    wire [64:0] _2815;
    wire [64:0] _2814;
    wire _2816;
    wire [63:0] _4904;
    wire [64:0] _2811;
    wire [64:0] _2802;
    wire [64:0] _2783;
    wire [64:0] _2782;
    wire _2784;
    wire [63:0] _4892;
    wire [64:0] _2779;
    wire [64:0] _2770;
    wire [64:0] _2751;
    wire [64:0] _2750;
    wire _2752;
    wire [63:0] _4880;
    wire [64:0] _2747;
    wire [64:0] _2738;
    wire [64:0] _2719;
    wire [64:0] _2718;
    wire _2720;
    wire [63:0] _4868;
    wire [64:0] _2715;
    wire [64:0] _2706;
    wire [64:0] _2687;
    wire [64:0] _2686;
    wire _2688;
    wire [63:0] _4856;
    wire [64:0] _2683;
    wire [64:0] _2674;
    wire [64:0] _2655;
    wire [64:0] _2654;
    wire _2656;
    wire [63:0] _4844;
    wire [64:0] _2651;
    wire [64:0] _2642;
    wire [64:0] _2623;
    wire [64:0] _2622;
    wire _2624;
    wire [63:0] _4832;
    wire [64:0] _2619;
    wire [64:0] _2610;
    wire [64:0] _2591;
    wire [64:0] _2590;
    wire _2592;
    wire [63:0] _4820;
    wire [64:0] _2587;
    wire [64:0] _2578;
    wire [64:0] _2559;
    wire [64:0] _2558;
    wire _2560;
    wire [63:0] _4808;
    wire [64:0] _2555;
    wire [64:0] _2546;
    wire [64:0] _2527;
    wire [64:0] _2526;
    wire _2528;
    wire [63:0] _4796;
    wire [64:0] _2523;
    wire [64:0] _2514;
    wire [64:0] _2495;
    wire [64:0] _2494;
    wire _2496;
    wire [63:0] _4784;
    wire [64:0] _2491;
    wire [64:0] _2482;
    wire [64:0] _2463;
    wire [64:0] _2462;
    wire _2464;
    wire [63:0] _4772;
    wire [64:0] _2459;
    wire [64:0] _2450;
    wire [64:0] _2431;
    wire [64:0] _2430;
    wire _2432;
    wire [63:0] _4760;
    wire [64:0] _2427;
    wire [64:0] _2418;
    wire [64:0] _2399;
    wire [64:0] _2398;
    wire _2400;
    wire [63:0] _4748;
    wire [64:0] _2395;
    wire [64:0] _2386;
    wire [64:0] _2367;
    wire [64:0] _2366;
    wire _2368;
    wire [63:0] _4736;
    wire [64:0] _2363;
    wire [64:0] _2354;
    wire [64:0] _2335;
    wire [64:0] _2334;
    wire _2336;
    wire [63:0] _4724;
    wire [64:0] _2331;
    wire [64:0] _2322;
    wire [64:0] _2303;
    wire [64:0] _2302;
    wire _2304;
    wire [63:0] _4712;
    wire [64:0] _2299;
    wire [64:0] _2290;
    wire [64:0] _2271;
    wire [64:0] _2270;
    wire _2272;
    wire [63:0] _4700;
    wire [64:0] _2267;
    wire [64:0] _2258;
    wire [64:0] _2239;
    wire [64:0] _2238;
    wire _2240;
    wire [63:0] _4688;
    wire [64:0] _2235;
    wire [64:0] _2226;
    wire [64:0] _2207;
    wire [64:0] _2206;
    wire _2208;
    wire [63:0] _4676;
    wire [64:0] _2203;
    wire [64:0] _2194;
    wire [64:0] _2175;
    wire [64:0] _2174;
    wire _2176;
    wire [63:0] _4664;
    wire [64:0] _2171;
    wire [64:0] _2162;
    wire [64:0] _2143;
    wire [64:0] _2142;
    wire _2144;
    wire [63:0] _4652;
    wire [64:0] _2139;
    wire [64:0] _2130;
    wire [64:0] _2111;
    wire [64:0] _2110;
    wire _2112;
    wire [63:0] _4640;
    wire [64:0] _2107;
    wire [64:0] _2098;
    wire [64:0] _2079;
    wire [64:0] _2078;
    wire _2080;
    wire [63:0] _4628;
    wire [64:0] _2075;
    wire [64:0] _2066;
    wire [64:0] _2047;
    wire [64:0] _2046;
    wire _2048;
    wire [63:0] _4616;
    wire [64:0] _2043;
    wire [64:0] _2034;
    wire [64:0] _2015;
    wire [64:0] _2014;
    wire _2016;
    wire [63:0] _4604;
    wire [64:0] _2011;
    wire [64:0] _2002;
    wire [64:0] _1983;
    wire [64:0] _1982;
    wire _1984;
    wire [63:0] _4592;
    wire [64:0] _1979;
    wire [64:0] _1970;
    wire [64:0] _1951;
    wire [64:0] _1950;
    wire _1952;
    wire [63:0] _4580;
    wire [64:0] _1947;
    wire [64:0] _1938;
    wire [64:0] _1919;
    wire [64:0] _1918;
    wire _1920;
    wire [63:0] _4568;
    wire [64:0] _1915;
    wire [64:0] _1906;
    wire [64:0] _1887;
    wire [64:0] _1886;
    wire _1888;
    wire [63:0] _4556;
    wire [64:0] _1883;
    wire [64:0] _1874;
    wire [64:0] _1855;
    wire [64:0] _1854;
    wire _1856;
    wire [63:0] _4544;
    wire [64:0] _1851;
    wire [64:0] _1842;
    wire [64:0] _1823;
    wire [64:0] _1822;
    wire _1824;
    wire [63:0] _4532;
    wire [64:0] _1819;
    wire [64:0] _1810;
    wire [64:0] _1791;
    wire [64:0] _1790;
    wire _1792;
    wire [63:0] _4520;
    wire [64:0] _1787;
    wire [64:0] _1778;
    wire [64:0] _1759;
    wire [64:0] _1758;
    wire _1760;
    wire [63:0] _4508;
    wire [64:0] _1755;
    wire [64:0] _1746;
    wire [64:0] _1727;
    wire [64:0] _1726;
    wire _1728;
    wire [63:0] _4496;
    wire [64:0] _1723;
    wire [64:0] _1714;
    wire [64:0] _1695;
    wire [64:0] _1694;
    wire _1696;
    wire [63:0] _4484;
    wire [64:0] _1691;
    wire [64:0] _1682;
    wire [64:0] _1663;
    wire [64:0] _1662;
    wire _1664;
    wire [63:0] _4472;
    wire [64:0] _1659;
    wire [64:0] _1650;
    wire [64:0] _1631;
    wire [64:0] _1630;
    wire _1632;
    wire [63:0] _4460;
    wire [64:0] _1627;
    wire [64:0] _1618;
    wire [64:0] _1599;
    wire [64:0] _1598;
    wire _1600;
    wire [63:0] _4448;
    wire [64:0] _1595;
    wire [64:0] _1586;
    wire [64:0] _1567;
    wire [64:0] _1566;
    wire _1568;
    wire [63:0] _4436;
    wire [64:0] _1563;
    wire [64:0] _1554;
    wire [64:0] _1535;
    wire [64:0] _1534;
    wire _1536;
    wire [63:0] _4424;
    wire [64:0] _1531;
    wire [64:0] _1522;
    wire [64:0] _1503;
    wire [64:0] _1502;
    wire _1504;
    wire [63:0] _4412;
    wire [64:0] _1499;
    wire [64:0] _1490;
    wire [64:0] _1471;
    wire [64:0] _1470;
    wire _1472;
    wire [63:0] _4400;
    wire [64:0] _1467;
    wire [64:0] _1458;
    wire [64:0] _1439;
    wire [64:0] _1438;
    wire _1440;
    wire [63:0] _4388;
    wire [64:0] _1435;
    wire [64:0] _1426;
    wire [64:0] _1407;
    wire [64:0] _1406;
    wire _1408;
    wire [63:0] _4376;
    wire [64:0] _1403;
    wire [64:0] _1394;
    wire [64:0] _1375;
    wire [64:0] _1374;
    wire _1376;
    wire [63:0] _4364;
    wire [64:0] _1371;
    wire [64:0] _1362;
    wire [64:0] _1343;
    wire [64:0] _1342;
    wire _1344;
    wire [63:0] _4352;
    wire [64:0] _1339;
    wire [64:0] _1330;
    wire [64:0] _1311;
    wire [64:0] _1310;
    wire _1312;
    wire [63:0] _4340;
    wire [64:0] _1307;
    wire [64:0] _1298;
    wire [64:0] _1279;
    wire [64:0] _1278;
    wire _1280;
    wire [63:0] _4328;
    wire [64:0] _1275;
    wire [64:0] _1266;
    wire [64:0] _1247;
    wire [64:0] _1246;
    wire _1248;
    wire [63:0] _4316;
    wire [64:0] _1243;
    wire [64:0] _1234;
    wire [64:0] _1215;
    wire [64:0] _1214;
    wire _1216;
    wire [63:0] _4304;
    wire [64:0] _1211;
    wire [64:0] _1202;
    wire [64:0] _1183;
    wire [64:0] _1182;
    wire _1184;
    wire [63:0] _4292;
    wire [64:0] _1179;
    wire [64:0] _1170;
    wire [64:0] _1151;
    wire [64:0] _1150;
    wire _1152;
    wire [63:0] _4280;
    wire [64:0] _1147;
    wire [64:0] _1138;
    wire [64:0] _1119;
    wire [64:0] _1118;
    wire _1120;
    wire [63:0] _4268;
    wire [64:0] _1115;
    wire [64:0] _1106;
    wire [64:0] _1087;
    wire [64:0] _1086;
    wire _1088;
    wire [63:0] _4256;
    wire [64:0] _1083;
    wire [64:0] _1074;
    wire [64:0] _1073;
    wire _1075;
    wire [63:0] _4250;
    wire [64:0] _1067;
    wire [64:0] _1066;
    wire _1068;
    wire [63:0] _4249;
    wire _1065;
    wire [63:0] _4251;
    wire [63:0] _4252;
    wire _4248;
    wire [63:0] _4253;
    wire [63:0] _205;
    reg [63:0] _1046;
    wire [64:0] _1082;
    wire _1084;
    wire [63:0] _4255;
    wire _1081;
    wire [63:0] _4257;
    wire [63:0] _4258;
    wire _4254;
    wire [63:0] _4259;
    wire [63:0] _206;
    reg [63:0] _1043;
    wire [64:0] _1105;
    wire _1107;
    wire [63:0] _4262;
    wire [64:0] _1099;
    wire [64:0] _1098;
    wire _1100;
    wire [63:0] _4261;
    wire _1097;
    wire [63:0] _4263;
    wire [63:0] _4264;
    wire _4260;
    wire [63:0] _4265;
    wire [63:0] _207;
    reg [63:0] _1040;
    wire [64:0] _1114;
    wire _1116;
    wire [63:0] _4267;
    wire _1113;
    wire [63:0] _4269;
    wire [63:0] _4270;
    wire _4266;
    wire [63:0] _4271;
    wire [63:0] _208;
    reg [63:0] _1037;
    wire [64:0] _1137;
    wire _1139;
    wire [63:0] _4274;
    wire [64:0] _1131;
    wire [64:0] _1130;
    wire _1132;
    wire [63:0] _4273;
    wire _1129;
    wire [63:0] _4275;
    wire [63:0] _4276;
    wire _4272;
    wire [63:0] _4277;
    wire [63:0] _209;
    reg [63:0] _1034;
    wire [64:0] _1146;
    wire _1148;
    wire [63:0] _4279;
    wire _1145;
    wire [63:0] _4281;
    wire [63:0] _4282;
    wire _4278;
    wire [63:0] _4283;
    wire [63:0] _210;
    reg [63:0] _1031;
    wire [64:0] _1169;
    wire _1171;
    wire [63:0] _4286;
    wire [64:0] _1163;
    wire [64:0] _1162;
    wire _1164;
    wire [63:0] _4285;
    wire _1161;
    wire [63:0] _4287;
    wire [63:0] _4288;
    wire _4284;
    wire [63:0] _4289;
    wire [63:0] _211;
    reg [63:0] _1028;
    wire [64:0] _1178;
    wire _1180;
    wire [63:0] _4291;
    wire _1177;
    wire [63:0] _4293;
    wire [63:0] _4294;
    wire _4290;
    wire [63:0] _4295;
    wire [63:0] _212;
    reg [63:0] _1025;
    wire [64:0] _1201;
    wire _1203;
    wire [63:0] _4298;
    wire [64:0] _1195;
    wire [64:0] _1194;
    wire _1196;
    wire [63:0] _4297;
    wire _1193;
    wire [63:0] _4299;
    wire [63:0] _4300;
    wire _4296;
    wire [63:0] _4301;
    wire [63:0] _213;
    reg [63:0] _1022;
    wire [64:0] _1210;
    wire _1212;
    wire [63:0] _4303;
    wire _1209;
    wire [63:0] _4305;
    wire [63:0] _4306;
    wire _4302;
    wire [63:0] _4307;
    wire [63:0] _214;
    reg [63:0] _1019;
    wire [64:0] _1233;
    wire _1235;
    wire [63:0] _4310;
    wire [64:0] _1227;
    wire [64:0] _1226;
    wire _1228;
    wire [63:0] _4309;
    wire _1225;
    wire [63:0] _4311;
    wire [63:0] _4312;
    wire _4308;
    wire [63:0] _4313;
    wire [63:0] _215;
    reg [63:0] _1016;
    wire [64:0] _1242;
    wire _1244;
    wire [63:0] _4315;
    wire _1241;
    wire [63:0] _4317;
    wire [63:0] _4318;
    wire _4314;
    wire [63:0] _4319;
    wire [63:0] _216;
    reg [63:0] _1013;
    wire [64:0] _1265;
    wire _1267;
    wire [63:0] _4322;
    wire [64:0] _1259;
    wire [64:0] _1258;
    wire _1260;
    wire [63:0] _4321;
    wire _1257;
    wire [63:0] _4323;
    wire [63:0] _4324;
    wire _4320;
    wire [63:0] _4325;
    wire [63:0] _217;
    reg [63:0] _1010;
    wire [64:0] _1274;
    wire _1276;
    wire [63:0] _4327;
    wire _1273;
    wire [63:0] _4329;
    wire [63:0] _4330;
    wire _4326;
    wire [63:0] _4331;
    wire [63:0] _218;
    reg [63:0] _1007;
    wire [64:0] _1297;
    wire _1299;
    wire [63:0] _4334;
    wire [64:0] _1291;
    wire [64:0] _1290;
    wire _1292;
    wire [63:0] _4333;
    wire _1289;
    wire [63:0] _4335;
    wire [63:0] _4336;
    wire _4332;
    wire [63:0] _4337;
    wire [63:0] _219;
    reg [63:0] _1004;
    wire [64:0] _1306;
    wire _1308;
    wire [63:0] _4339;
    wire _1305;
    wire [63:0] _4341;
    wire [63:0] _4342;
    wire _4338;
    wire [63:0] _4343;
    wire [63:0] _220;
    reg [63:0] _1001;
    wire [64:0] _1329;
    wire _1331;
    wire [63:0] _4346;
    wire [64:0] _1323;
    wire [64:0] _1322;
    wire _1324;
    wire [63:0] _4345;
    wire _1321;
    wire [63:0] _4347;
    wire [63:0] _4348;
    wire _4344;
    wire [63:0] _4349;
    wire [63:0] _221;
    reg [63:0] _998;
    wire [64:0] _1338;
    wire _1340;
    wire [63:0] _4351;
    wire _1337;
    wire [63:0] _4353;
    wire [63:0] _4354;
    wire _4350;
    wire [63:0] _4355;
    wire [63:0] _222;
    reg [63:0] _995;
    wire [64:0] _1361;
    wire _1363;
    wire [63:0] _4358;
    wire [64:0] _1355;
    wire [64:0] _1354;
    wire _1356;
    wire [63:0] _4357;
    wire _1353;
    wire [63:0] _4359;
    wire [63:0] _4360;
    wire _4356;
    wire [63:0] _4361;
    wire [63:0] _223;
    reg [63:0] _992;
    wire [64:0] _1370;
    wire _1372;
    wire [63:0] _4363;
    wire _1369;
    wire [63:0] _4365;
    wire [63:0] _4366;
    wire _4362;
    wire [63:0] _4367;
    wire [63:0] _224;
    reg [63:0] _989;
    wire [64:0] _1393;
    wire _1395;
    wire [63:0] _4370;
    wire [64:0] _1387;
    wire [64:0] _1386;
    wire _1388;
    wire [63:0] _4369;
    wire _1385;
    wire [63:0] _4371;
    wire [63:0] _4372;
    wire _4368;
    wire [63:0] _4373;
    wire [63:0] _225;
    reg [63:0] _986;
    wire [64:0] _1402;
    wire _1404;
    wire [63:0] _4375;
    wire _1401;
    wire [63:0] _4377;
    wire [63:0] _4378;
    wire _4374;
    wire [63:0] _4379;
    wire [63:0] _226;
    reg [63:0] _983;
    wire [64:0] _1425;
    wire _1427;
    wire [63:0] _4382;
    wire [64:0] _1419;
    wire [64:0] _1418;
    wire _1420;
    wire [63:0] _4381;
    wire _1417;
    wire [63:0] _4383;
    wire [63:0] _4384;
    wire _4380;
    wire [63:0] _4385;
    wire [63:0] _227;
    reg [63:0] _980;
    wire [64:0] _1434;
    wire _1436;
    wire [63:0] _4387;
    wire _1433;
    wire [63:0] _4389;
    wire [63:0] _4390;
    wire _4386;
    wire [63:0] _4391;
    wire [63:0] _228;
    reg [63:0] _977;
    wire [64:0] _1457;
    wire _1459;
    wire [63:0] _4394;
    wire [64:0] _1451;
    wire [64:0] _1450;
    wire _1452;
    wire [63:0] _4393;
    wire _1449;
    wire [63:0] _4395;
    wire [63:0] _4396;
    wire _4392;
    wire [63:0] _4397;
    wire [63:0] _229;
    reg [63:0] _974;
    wire [64:0] _1466;
    wire _1468;
    wire [63:0] _4399;
    wire _1465;
    wire [63:0] _4401;
    wire [63:0] _4402;
    wire _4398;
    wire [63:0] _4403;
    wire [63:0] _230;
    reg [63:0] _971;
    wire [64:0] _1489;
    wire _1491;
    wire [63:0] _4406;
    wire [64:0] _1483;
    wire [64:0] _1482;
    wire _1484;
    wire [63:0] _4405;
    wire _1481;
    wire [63:0] _4407;
    wire [63:0] _4408;
    wire _4404;
    wire [63:0] _4409;
    wire [63:0] _231;
    reg [63:0] _968;
    wire [64:0] _1498;
    wire _1500;
    wire [63:0] _4411;
    wire _1497;
    wire [63:0] _4413;
    wire [63:0] _4414;
    wire _4410;
    wire [63:0] _4415;
    wire [63:0] _232;
    reg [63:0] _965;
    wire [64:0] _1521;
    wire _1523;
    wire [63:0] _4418;
    wire [64:0] _1515;
    wire [64:0] _1514;
    wire _1516;
    wire [63:0] _4417;
    wire _1513;
    wire [63:0] _4419;
    wire [63:0] _4420;
    wire _4416;
    wire [63:0] _4421;
    wire [63:0] _233;
    reg [63:0] _962;
    wire [64:0] _1530;
    wire _1532;
    wire [63:0] _4423;
    wire _1529;
    wire [63:0] _4425;
    wire [63:0] _4426;
    wire _4422;
    wire [63:0] _4427;
    wire [63:0] _234;
    reg [63:0] _959;
    wire [64:0] _1553;
    wire _1555;
    wire [63:0] _4430;
    wire [64:0] _1547;
    wire [64:0] _1546;
    wire _1548;
    wire [63:0] _4429;
    wire _1545;
    wire [63:0] _4431;
    wire [63:0] _4432;
    wire _4428;
    wire [63:0] _4433;
    wire [63:0] _235;
    reg [63:0] _956;
    wire [64:0] _1562;
    wire _1564;
    wire [63:0] _4435;
    wire _1561;
    wire [63:0] _4437;
    wire [63:0] _4438;
    wire _4434;
    wire [63:0] _4439;
    wire [63:0] _236;
    reg [63:0] _953;
    wire [64:0] _1585;
    wire _1587;
    wire [63:0] _4442;
    wire [64:0] _1579;
    wire [64:0] _1578;
    wire _1580;
    wire [63:0] _4441;
    wire _1577;
    wire [63:0] _4443;
    wire [63:0] _4444;
    wire _4440;
    wire [63:0] _4445;
    wire [63:0] _237;
    reg [63:0] _950;
    wire [64:0] _1594;
    wire _1596;
    wire [63:0] _4447;
    wire _1593;
    wire [63:0] _4449;
    wire [63:0] _4450;
    wire _4446;
    wire [63:0] _4451;
    wire [63:0] _238;
    reg [63:0] _947;
    wire [64:0] _1617;
    wire _1619;
    wire [63:0] _4454;
    wire [64:0] _1611;
    wire [64:0] _1610;
    wire _1612;
    wire [63:0] _4453;
    wire _1609;
    wire [63:0] _4455;
    wire [63:0] _4456;
    wire _4452;
    wire [63:0] _4457;
    wire [63:0] _239;
    reg [63:0] _944;
    wire [64:0] _1626;
    wire _1628;
    wire [63:0] _4459;
    wire _1625;
    wire [63:0] _4461;
    wire [63:0] _4462;
    wire _4458;
    wire [63:0] _4463;
    wire [63:0] _240;
    reg [63:0] _941;
    wire [64:0] _1649;
    wire _1651;
    wire [63:0] _4466;
    wire [64:0] _1643;
    wire [64:0] _1642;
    wire _1644;
    wire [63:0] _4465;
    wire _1641;
    wire [63:0] _4467;
    wire [63:0] _4468;
    wire _4464;
    wire [63:0] _4469;
    wire [63:0] _241;
    reg [63:0] _938;
    wire [64:0] _1658;
    wire _1660;
    wire [63:0] _4471;
    wire _1657;
    wire [63:0] _4473;
    wire [63:0] _4474;
    wire _4470;
    wire [63:0] _4475;
    wire [63:0] _242;
    reg [63:0] _935;
    wire [64:0] _1681;
    wire _1683;
    wire [63:0] _4478;
    wire [64:0] _1675;
    wire [64:0] _1674;
    wire _1676;
    wire [63:0] _4477;
    wire _1673;
    wire [63:0] _4479;
    wire [63:0] _4480;
    wire _4476;
    wire [63:0] _4481;
    wire [63:0] _243;
    reg [63:0] _932;
    wire [64:0] _1690;
    wire _1692;
    wire [63:0] _4483;
    wire _1689;
    wire [63:0] _4485;
    wire [63:0] _4486;
    wire _4482;
    wire [63:0] _4487;
    wire [63:0] _244;
    reg [63:0] _929;
    wire [64:0] _1713;
    wire _1715;
    wire [63:0] _4490;
    wire [64:0] _1707;
    wire [64:0] _1706;
    wire _1708;
    wire [63:0] _4489;
    wire _1705;
    wire [63:0] _4491;
    wire [63:0] _4492;
    wire _4488;
    wire [63:0] _4493;
    wire [63:0] _245;
    reg [63:0] _926;
    wire [64:0] _1722;
    wire _1724;
    wire [63:0] _4495;
    wire _1721;
    wire [63:0] _4497;
    wire [63:0] _4498;
    wire _4494;
    wire [63:0] _4499;
    wire [63:0] _246;
    reg [63:0] _923;
    wire [64:0] _1745;
    wire _1747;
    wire [63:0] _4502;
    wire [64:0] _1739;
    wire [64:0] _1738;
    wire _1740;
    wire [63:0] _4501;
    wire _1737;
    wire [63:0] _4503;
    wire [63:0] _4504;
    wire _4500;
    wire [63:0] _4505;
    wire [63:0] _247;
    reg [63:0] _920;
    wire [64:0] _1754;
    wire _1756;
    wire [63:0] _4507;
    wire _1753;
    wire [63:0] _4509;
    wire [63:0] _4510;
    wire _4506;
    wire [63:0] _4511;
    wire [63:0] _248;
    reg [63:0] _917;
    wire [64:0] _1777;
    wire _1779;
    wire [63:0] _4514;
    wire [64:0] _1771;
    wire [64:0] _1770;
    wire _1772;
    wire [63:0] _4513;
    wire _1769;
    wire [63:0] _4515;
    wire [63:0] _4516;
    wire _4512;
    wire [63:0] _4517;
    wire [63:0] _249;
    reg [63:0] _914;
    wire [64:0] _1786;
    wire _1788;
    wire [63:0] _4519;
    wire _1785;
    wire [63:0] _4521;
    wire [63:0] _4522;
    wire _4518;
    wire [63:0] _4523;
    wire [63:0] _250;
    reg [63:0] _911;
    wire [64:0] _1809;
    wire _1811;
    wire [63:0] _4526;
    wire [64:0] _1803;
    wire [64:0] _1802;
    wire _1804;
    wire [63:0] _4525;
    wire _1801;
    wire [63:0] _4527;
    wire [63:0] _4528;
    wire _4524;
    wire [63:0] _4529;
    wire [63:0] _251;
    reg [63:0] _908;
    wire [64:0] _1818;
    wire _1820;
    wire [63:0] _4531;
    wire _1817;
    wire [63:0] _4533;
    wire [63:0] _4534;
    wire _4530;
    wire [63:0] _4535;
    wire [63:0] _252;
    reg [63:0] _905;
    wire [64:0] _1841;
    wire _1843;
    wire [63:0] _4538;
    wire [64:0] _1835;
    wire [64:0] _1834;
    wire _1836;
    wire [63:0] _4537;
    wire _1833;
    wire [63:0] _4539;
    wire [63:0] _4540;
    wire _4536;
    wire [63:0] _4541;
    wire [63:0] _253;
    reg [63:0] _902;
    wire [64:0] _1850;
    wire _1852;
    wire [63:0] _4543;
    wire _1849;
    wire [63:0] _4545;
    wire [63:0] _4546;
    wire _4542;
    wire [63:0] _4547;
    wire [63:0] _254;
    reg [63:0] _899;
    wire [64:0] _1873;
    wire _1875;
    wire [63:0] _4550;
    wire [64:0] _1867;
    wire [64:0] _1866;
    wire _1868;
    wire [63:0] _4549;
    wire _1865;
    wire [63:0] _4551;
    wire [63:0] _4552;
    wire _4548;
    wire [63:0] _4553;
    wire [63:0] _255;
    reg [63:0] _896;
    wire [64:0] _1882;
    wire _1884;
    wire [63:0] _4555;
    wire _1881;
    wire [63:0] _4557;
    wire [63:0] _4558;
    wire _4554;
    wire [63:0] _4559;
    wire [63:0] _256;
    reg [63:0] _893;
    wire [64:0] _1905;
    wire _1907;
    wire [63:0] _4562;
    wire [64:0] _1899;
    wire [64:0] _1898;
    wire _1900;
    wire [63:0] _4561;
    wire _1897;
    wire [63:0] _4563;
    wire [63:0] _4564;
    wire _4560;
    wire [63:0] _4565;
    wire [63:0] _257;
    reg [63:0] _890;
    wire [64:0] _1914;
    wire _1916;
    wire [63:0] _4567;
    wire _1913;
    wire [63:0] _4569;
    wire [63:0] _4570;
    wire _4566;
    wire [63:0] _4571;
    wire [63:0] _258;
    reg [63:0] _887;
    wire [64:0] _1937;
    wire _1939;
    wire [63:0] _4574;
    wire [64:0] _1931;
    wire [64:0] _1930;
    wire _1932;
    wire [63:0] _4573;
    wire _1929;
    wire [63:0] _4575;
    wire [63:0] _4576;
    wire _4572;
    wire [63:0] _4577;
    wire [63:0] _259;
    reg [63:0] _884;
    wire [64:0] _1946;
    wire _1948;
    wire [63:0] _4579;
    wire _1945;
    wire [63:0] _4581;
    wire [63:0] _4582;
    wire _4578;
    wire [63:0] _4583;
    wire [63:0] _260;
    reg [63:0] _881;
    wire [64:0] _1969;
    wire _1971;
    wire [63:0] _4586;
    wire [64:0] _1963;
    wire [64:0] _1962;
    wire _1964;
    wire [63:0] _4585;
    wire _1961;
    wire [63:0] _4587;
    wire [63:0] _4588;
    wire _4584;
    wire [63:0] _4589;
    wire [63:0] _261;
    reg [63:0] _878;
    wire [64:0] _1978;
    wire _1980;
    wire [63:0] _4591;
    wire _1977;
    wire [63:0] _4593;
    wire [63:0] _4594;
    wire _4590;
    wire [63:0] _4595;
    wire [63:0] _262;
    reg [63:0] _875;
    wire [64:0] _2001;
    wire _2003;
    wire [63:0] _4598;
    wire [64:0] _1995;
    wire [64:0] _1994;
    wire _1996;
    wire [63:0] _4597;
    wire _1993;
    wire [63:0] _4599;
    wire [63:0] _4600;
    wire _4596;
    wire [63:0] _4601;
    wire [63:0] _263;
    reg [63:0] _872;
    wire [64:0] _2010;
    wire _2012;
    wire [63:0] _4603;
    wire _2009;
    wire [63:0] _4605;
    wire [63:0] _4606;
    wire _4602;
    wire [63:0] _4607;
    wire [63:0] _264;
    reg [63:0] _869;
    wire [64:0] _2033;
    wire _2035;
    wire [63:0] _4610;
    wire [64:0] _2027;
    wire [64:0] _2026;
    wire _2028;
    wire [63:0] _4609;
    wire _2025;
    wire [63:0] _4611;
    wire [63:0] _4612;
    wire _4608;
    wire [63:0] _4613;
    wire [63:0] _265;
    reg [63:0] _866;
    wire [64:0] _2042;
    wire _2044;
    wire [63:0] _4615;
    wire _2041;
    wire [63:0] _4617;
    wire [63:0] _4618;
    wire _4614;
    wire [63:0] _4619;
    wire [63:0] _266;
    reg [63:0] _863;
    wire [64:0] _2065;
    wire _2067;
    wire [63:0] _4622;
    wire [64:0] _2059;
    wire [64:0] _2058;
    wire _2060;
    wire [63:0] _4621;
    wire _2057;
    wire [63:0] _4623;
    wire [63:0] _4624;
    wire _4620;
    wire [63:0] _4625;
    wire [63:0] _267;
    reg [63:0] _860;
    wire [64:0] _2074;
    wire _2076;
    wire [63:0] _4627;
    wire _2073;
    wire [63:0] _4629;
    wire [63:0] _4630;
    wire _4626;
    wire [63:0] _4631;
    wire [63:0] _268;
    reg [63:0] _857;
    wire [64:0] _2097;
    wire _2099;
    wire [63:0] _4634;
    wire [64:0] _2091;
    wire [64:0] _2090;
    wire _2092;
    wire [63:0] _4633;
    wire _2089;
    wire [63:0] _4635;
    wire [63:0] _4636;
    wire _4632;
    wire [63:0] _4637;
    wire [63:0] _269;
    reg [63:0] _854;
    wire [64:0] _2106;
    wire _2108;
    wire [63:0] _4639;
    wire _2105;
    wire [63:0] _4641;
    wire [63:0] _4642;
    wire _4638;
    wire [63:0] _4643;
    wire [63:0] _270;
    reg [63:0] _851;
    wire [64:0] _2129;
    wire _2131;
    wire [63:0] _4646;
    wire [64:0] _2123;
    wire [64:0] _2122;
    wire _2124;
    wire [63:0] _4645;
    wire _2121;
    wire [63:0] _4647;
    wire [63:0] _4648;
    wire _4644;
    wire [63:0] _4649;
    wire [63:0] _271;
    reg [63:0] _848;
    wire [64:0] _2138;
    wire _2140;
    wire [63:0] _4651;
    wire _2137;
    wire [63:0] _4653;
    wire [63:0] _4654;
    wire _4650;
    wire [63:0] _4655;
    wire [63:0] _272;
    reg [63:0] _845;
    wire [64:0] _2161;
    wire _2163;
    wire [63:0] _4658;
    wire [64:0] _2155;
    wire [64:0] _2154;
    wire _2156;
    wire [63:0] _4657;
    wire _2153;
    wire [63:0] _4659;
    wire [63:0] _4660;
    wire _4656;
    wire [63:0] _4661;
    wire [63:0] _273;
    reg [63:0] _842;
    wire [64:0] _2170;
    wire _2172;
    wire [63:0] _4663;
    wire _2169;
    wire [63:0] _4665;
    wire [63:0] _4666;
    wire _4662;
    wire [63:0] _4667;
    wire [63:0] _274;
    reg [63:0] _839;
    wire [64:0] _2193;
    wire _2195;
    wire [63:0] _4670;
    wire [64:0] _2187;
    wire [64:0] _2186;
    wire _2188;
    wire [63:0] _4669;
    wire _2185;
    wire [63:0] _4671;
    wire [63:0] _4672;
    wire _4668;
    wire [63:0] _4673;
    wire [63:0] _275;
    reg [63:0] _836;
    wire [64:0] _2202;
    wire _2204;
    wire [63:0] _4675;
    wire _2201;
    wire [63:0] _4677;
    wire [63:0] _4678;
    wire _4674;
    wire [63:0] _4679;
    wire [63:0] _276;
    reg [63:0] _833;
    wire [64:0] _2225;
    wire _2227;
    wire [63:0] _4682;
    wire [64:0] _2219;
    wire [64:0] _2218;
    wire _2220;
    wire [63:0] _4681;
    wire _2217;
    wire [63:0] _4683;
    wire [63:0] _4684;
    wire _4680;
    wire [63:0] _4685;
    wire [63:0] _277;
    reg [63:0] _830;
    wire [64:0] _2234;
    wire _2236;
    wire [63:0] _4687;
    wire _2233;
    wire [63:0] _4689;
    wire [63:0] _4690;
    wire _4686;
    wire [63:0] _4691;
    wire [63:0] _278;
    reg [63:0] _827;
    wire [64:0] _2257;
    wire _2259;
    wire [63:0] _4694;
    wire [64:0] _2251;
    wire [64:0] _2250;
    wire _2252;
    wire [63:0] _4693;
    wire _2249;
    wire [63:0] _4695;
    wire [63:0] _4696;
    wire _4692;
    wire [63:0] _4697;
    wire [63:0] _279;
    reg [63:0] _824;
    wire [64:0] _2266;
    wire _2268;
    wire [63:0] _4699;
    wire _2265;
    wire [63:0] _4701;
    wire [63:0] _4702;
    wire _4698;
    wire [63:0] _4703;
    wire [63:0] _280;
    reg [63:0] _821;
    wire [64:0] _2289;
    wire _2291;
    wire [63:0] _4706;
    wire [64:0] _2283;
    wire [64:0] _2282;
    wire _2284;
    wire [63:0] _4705;
    wire _2281;
    wire [63:0] _4707;
    wire [63:0] _4708;
    wire _4704;
    wire [63:0] _4709;
    wire [63:0] _281;
    reg [63:0] _818;
    wire [64:0] _2298;
    wire _2300;
    wire [63:0] _4711;
    wire _2297;
    wire [63:0] _4713;
    wire [63:0] _4714;
    wire _4710;
    wire [63:0] _4715;
    wire [63:0] _282;
    reg [63:0] _815;
    wire [64:0] _2321;
    wire _2323;
    wire [63:0] _4718;
    wire [64:0] _2315;
    wire [64:0] _2314;
    wire _2316;
    wire [63:0] _4717;
    wire _2313;
    wire [63:0] _4719;
    wire [63:0] _4720;
    wire _4716;
    wire [63:0] _4721;
    wire [63:0] _283;
    reg [63:0] _812;
    wire [64:0] _2330;
    wire _2332;
    wire [63:0] _4723;
    wire _2329;
    wire [63:0] _4725;
    wire [63:0] _4726;
    wire _4722;
    wire [63:0] _4727;
    wire [63:0] _284;
    reg [63:0] _809;
    wire [64:0] _2353;
    wire _2355;
    wire [63:0] _4730;
    wire [64:0] _2347;
    wire [64:0] _2346;
    wire _2348;
    wire [63:0] _4729;
    wire _2345;
    wire [63:0] _4731;
    wire [63:0] _4732;
    wire _4728;
    wire [63:0] _4733;
    wire [63:0] _285;
    reg [63:0] _806;
    wire [64:0] _2362;
    wire _2364;
    wire [63:0] _4735;
    wire _2361;
    wire [63:0] _4737;
    wire [63:0] _4738;
    wire _4734;
    wire [63:0] _4739;
    wire [63:0] _286;
    reg [63:0] _803;
    wire [64:0] _2385;
    wire _2387;
    wire [63:0] _4742;
    wire [64:0] _2379;
    wire [64:0] _2378;
    wire _2380;
    wire [63:0] _4741;
    wire _2377;
    wire [63:0] _4743;
    wire [63:0] _4744;
    wire _4740;
    wire [63:0] _4745;
    wire [63:0] _287;
    reg [63:0] _800;
    wire [64:0] _2394;
    wire _2396;
    wire [63:0] _4747;
    wire _2393;
    wire [63:0] _4749;
    wire [63:0] _4750;
    wire _4746;
    wire [63:0] _4751;
    wire [63:0] _288;
    reg [63:0] _797;
    wire [64:0] _2417;
    wire _2419;
    wire [63:0] _4754;
    wire [64:0] _2411;
    wire [64:0] _2410;
    wire _2412;
    wire [63:0] _4753;
    wire _2409;
    wire [63:0] _4755;
    wire [63:0] _4756;
    wire _4752;
    wire [63:0] _4757;
    wire [63:0] _289;
    reg [63:0] _794;
    wire [64:0] _2426;
    wire _2428;
    wire [63:0] _4759;
    wire _2425;
    wire [63:0] _4761;
    wire [63:0] _4762;
    wire _4758;
    wire [63:0] _4763;
    wire [63:0] _290;
    reg [63:0] _791;
    wire [64:0] _2449;
    wire _2451;
    wire [63:0] _4766;
    wire [64:0] _2443;
    wire [64:0] _2442;
    wire _2444;
    wire [63:0] _4765;
    wire _2441;
    wire [63:0] _4767;
    wire [63:0] _4768;
    wire _4764;
    wire [63:0] _4769;
    wire [63:0] _291;
    reg [63:0] _788;
    wire [64:0] _2458;
    wire _2460;
    wire [63:0] _4771;
    wire _2457;
    wire [63:0] _4773;
    wire [63:0] _4774;
    wire _4770;
    wire [63:0] _4775;
    wire [63:0] _292;
    reg [63:0] _785;
    wire [64:0] _2481;
    wire _2483;
    wire [63:0] _4778;
    wire [64:0] _2475;
    wire [64:0] _2474;
    wire _2476;
    wire [63:0] _4777;
    wire _2473;
    wire [63:0] _4779;
    wire [63:0] _4780;
    wire _4776;
    wire [63:0] _4781;
    wire [63:0] _293;
    reg [63:0] _782;
    wire [64:0] _2490;
    wire _2492;
    wire [63:0] _4783;
    wire _2489;
    wire [63:0] _4785;
    wire [63:0] _4786;
    wire _4782;
    wire [63:0] _4787;
    wire [63:0] _294;
    reg [63:0] _779;
    wire [64:0] _2513;
    wire _2515;
    wire [63:0] _4790;
    wire [64:0] _2507;
    wire [64:0] _2506;
    wire _2508;
    wire [63:0] _4789;
    wire _2505;
    wire [63:0] _4791;
    wire [63:0] _4792;
    wire _4788;
    wire [63:0] _4793;
    wire [63:0] _295;
    reg [63:0] _776;
    wire [64:0] _2522;
    wire _2524;
    wire [63:0] _4795;
    wire _2521;
    wire [63:0] _4797;
    wire [63:0] _4798;
    wire _4794;
    wire [63:0] _4799;
    wire [63:0] _296;
    reg [63:0] _773;
    wire [64:0] _2545;
    wire _2547;
    wire [63:0] _4802;
    wire [64:0] _2539;
    wire [64:0] _2538;
    wire _2540;
    wire [63:0] _4801;
    wire _2537;
    wire [63:0] _4803;
    wire [63:0] _4804;
    wire _4800;
    wire [63:0] _4805;
    wire [63:0] _297;
    reg [63:0] _770;
    wire [64:0] _2554;
    wire _2556;
    wire [63:0] _4807;
    wire _2553;
    wire [63:0] _4809;
    wire [63:0] _4810;
    wire _4806;
    wire [63:0] _4811;
    wire [63:0] _298;
    reg [63:0] _767;
    wire [64:0] _2577;
    wire _2579;
    wire [63:0] _4814;
    wire [64:0] _2571;
    wire [64:0] _2570;
    wire _2572;
    wire [63:0] _4813;
    wire _2569;
    wire [63:0] _4815;
    wire [63:0] _4816;
    wire _4812;
    wire [63:0] _4817;
    wire [63:0] _299;
    reg [63:0] _764;
    wire [64:0] _2586;
    wire _2588;
    wire [63:0] _4819;
    wire _2585;
    wire [63:0] _4821;
    wire [63:0] _4822;
    wire _4818;
    wire [63:0] _4823;
    wire [63:0] _300;
    reg [63:0] _761;
    wire [64:0] _2609;
    wire _2611;
    wire [63:0] _4826;
    wire [64:0] _2603;
    wire [64:0] _2602;
    wire _2604;
    wire [63:0] _4825;
    wire _2601;
    wire [63:0] _4827;
    wire [63:0] _4828;
    wire _4824;
    wire [63:0] _4829;
    wire [63:0] _301;
    reg [63:0] _758;
    wire [64:0] _2618;
    wire _2620;
    wire [63:0] _4831;
    wire _2617;
    wire [63:0] _4833;
    wire [63:0] _4834;
    wire _4830;
    wire [63:0] _4835;
    wire [63:0] _302;
    reg [63:0] _755;
    wire [64:0] _2641;
    wire _2643;
    wire [63:0] _4838;
    wire [64:0] _2635;
    wire [64:0] _2634;
    wire _2636;
    wire [63:0] _4837;
    wire _2633;
    wire [63:0] _4839;
    wire [63:0] _4840;
    wire _4836;
    wire [63:0] _4841;
    wire [63:0] _303;
    reg [63:0] _752;
    wire [64:0] _2650;
    wire _2652;
    wire [63:0] _4843;
    wire _2649;
    wire [63:0] _4845;
    wire [63:0] _4846;
    wire _4842;
    wire [63:0] _4847;
    wire [63:0] _304;
    reg [63:0] _749;
    wire [64:0] _2673;
    wire _2675;
    wire [63:0] _4850;
    wire [64:0] _2667;
    wire [64:0] _2666;
    wire _2668;
    wire [63:0] _4849;
    wire _2665;
    wire [63:0] _4851;
    wire [63:0] _4852;
    wire _4848;
    wire [63:0] _4853;
    wire [63:0] _305;
    reg [63:0] _746;
    wire [64:0] _2682;
    wire _2684;
    wire [63:0] _4855;
    wire _2681;
    wire [63:0] _4857;
    wire [63:0] _4858;
    wire _4854;
    wire [63:0] _4859;
    wire [63:0] _306;
    reg [63:0] _743;
    wire [64:0] _2705;
    wire _2707;
    wire [63:0] _4862;
    wire [64:0] _2699;
    wire [64:0] _2698;
    wire _2700;
    wire [63:0] _4861;
    wire _2697;
    wire [63:0] _4863;
    wire [63:0] _4864;
    wire _4860;
    wire [63:0] _4865;
    wire [63:0] _307;
    reg [63:0] _740;
    wire [64:0] _2714;
    wire _2716;
    wire [63:0] _4867;
    wire _2713;
    wire [63:0] _4869;
    wire [63:0] _4870;
    wire _4866;
    wire [63:0] _4871;
    wire [63:0] _308;
    reg [63:0] _737;
    wire [64:0] _2737;
    wire _2739;
    wire [63:0] _4874;
    wire [64:0] _2731;
    wire [64:0] _2730;
    wire _2732;
    wire [63:0] _4873;
    wire _2729;
    wire [63:0] _4875;
    wire [63:0] _4876;
    wire _4872;
    wire [63:0] _4877;
    wire [63:0] _309;
    reg [63:0] _734;
    wire [64:0] _2746;
    wire _2748;
    wire [63:0] _4879;
    wire _2745;
    wire [63:0] _4881;
    wire [63:0] _4882;
    wire _4878;
    wire [63:0] _4883;
    wire [63:0] _310;
    reg [63:0] _731;
    wire [64:0] _2769;
    wire _2771;
    wire [63:0] _4886;
    wire [64:0] _2763;
    wire [64:0] _2762;
    wire _2764;
    wire [63:0] _4885;
    wire _2761;
    wire [63:0] _4887;
    wire [63:0] _4888;
    wire _4884;
    wire [63:0] _4889;
    wire [63:0] _311;
    reg [63:0] _728;
    wire [64:0] _2778;
    wire _2780;
    wire [63:0] _4891;
    wire _2777;
    wire [63:0] _4893;
    wire [63:0] _4894;
    wire _4890;
    wire [63:0] _4895;
    wire [63:0] _312;
    reg [63:0] _725;
    wire [64:0] _2801;
    wire _2803;
    wire [63:0] _4898;
    wire [64:0] _2795;
    wire [64:0] _2794;
    wire _2796;
    wire [63:0] _4897;
    wire _2793;
    wire [63:0] _4899;
    wire [63:0] _4900;
    wire _4896;
    wire [63:0] _4901;
    wire [63:0] _313;
    reg [63:0] _722;
    wire [64:0] _2810;
    wire _2812;
    wire [63:0] _4903;
    wire _2809;
    wire [63:0] _4905;
    wire [63:0] _4906;
    wire _4902;
    wire [63:0] _4907;
    wire [63:0] _314;
    reg [63:0] _719;
    wire [64:0] _2833;
    wire _2835;
    wire [63:0] _4910;
    wire [64:0] _2827;
    wire [64:0] _2826;
    wire _2828;
    wire [63:0] _4909;
    wire _2825;
    wire [63:0] _4911;
    wire [63:0] _4912;
    wire _4908;
    wire [63:0] _4913;
    wire [63:0] _315;
    reg [63:0] _716;
    wire [64:0] _2842;
    wire _2844;
    wire [63:0] _4915;
    wire _2841;
    wire [63:0] _4917;
    wire [63:0] _4918;
    wire _4914;
    wire [63:0] _4919;
    wire [63:0] _316;
    reg [63:0] _713;
    wire [64:0] _2865;
    wire _2867;
    wire [63:0] _4922;
    wire [64:0] _2859;
    wire [64:0] _2858;
    wire _2860;
    wire [63:0] _4921;
    wire _2857;
    wire [63:0] _4923;
    wire [63:0] _4924;
    wire _4920;
    wire [63:0] _4925;
    wire [63:0] _317;
    reg [63:0] _710;
    wire [64:0] _2874;
    wire _2876;
    wire [63:0] _4927;
    wire _2873;
    wire [63:0] _4929;
    wire [63:0] _4930;
    wire _4926;
    wire [63:0] _4931;
    wire [63:0] _318;
    reg [63:0] _707;
    wire [64:0] _2897;
    wire _2899;
    wire [63:0] _4934;
    wire [64:0] _2891;
    wire [64:0] _2890;
    wire _2892;
    wire [63:0] _4933;
    wire _2889;
    wire [63:0] _4935;
    wire [63:0] _4936;
    wire _4932;
    wire [63:0] _4937;
    wire [63:0] _319;
    reg [63:0] _704;
    wire [64:0] _2906;
    wire _2908;
    wire [63:0] _4939;
    wire _2905;
    wire [63:0] _4941;
    wire [63:0] _4942;
    wire _4938;
    wire [63:0] _4943;
    wire [63:0] _320;
    reg [63:0] _701;
    wire [64:0] _2929;
    wire _2931;
    wire [63:0] _4946;
    wire [64:0] _2923;
    wire [64:0] _2922;
    wire _2924;
    wire [63:0] _4945;
    wire _2921;
    wire [63:0] _4947;
    wire [63:0] _4948;
    wire _4944;
    wire [63:0] _4949;
    wire [63:0] _321;
    reg [63:0] _698;
    wire [64:0] _2938;
    wire _2940;
    wire [63:0] _4951;
    wire _2937;
    wire [63:0] _4953;
    wire [63:0] _4954;
    wire _4950;
    wire [63:0] _4955;
    wire [63:0] _322;
    reg [63:0] _695;
    wire [64:0] _2961;
    wire _2963;
    wire [63:0] _4958;
    wire [64:0] _2955;
    wire [64:0] _2954;
    wire _2956;
    wire [63:0] _4957;
    wire _2953;
    wire [63:0] _4959;
    wire [63:0] _4960;
    wire _4956;
    wire [63:0] _4961;
    wire [63:0] _323;
    reg [63:0] _692;
    wire [64:0] _2970;
    wire _2972;
    wire [63:0] _4963;
    wire _2969;
    wire [63:0] _4965;
    wire [63:0] _4966;
    wire _4962;
    wire [63:0] _4967;
    wire [63:0] _324;
    reg [63:0] _689;
    wire [64:0] _2993;
    wire _2995;
    wire [63:0] _4970;
    wire [64:0] _2987;
    wire [64:0] _2986;
    wire _2988;
    wire [63:0] _4969;
    wire _2985;
    wire [63:0] _4971;
    wire [63:0] _4972;
    wire _4968;
    wire [63:0] _4973;
    wire [63:0] _325;
    reg [63:0] _686;
    wire [64:0] _3002;
    wire _3004;
    wire [63:0] _4975;
    wire _3001;
    wire [63:0] _4977;
    wire [63:0] _4978;
    wire _4974;
    wire [63:0] _4979;
    wire [63:0] _326;
    reg [63:0] _683;
    wire [64:0] _3025;
    wire _3027;
    wire [63:0] _4982;
    wire [64:0] _3019;
    wire [64:0] _3018;
    wire _3020;
    wire [63:0] _4981;
    wire _3017;
    wire [63:0] _4983;
    wire [63:0] _4984;
    wire _4980;
    wire [63:0] _4985;
    wire [63:0] _327;
    reg [63:0] _680;
    wire [64:0] _3034;
    wire _3036;
    wire [63:0] _4987;
    wire _3033;
    wire [63:0] _4989;
    wire [63:0] _4990;
    wire _4986;
    wire [63:0] _4991;
    wire [63:0] _328;
    reg [63:0] _677;
    wire [64:0] _3057;
    wire _3059;
    wire [63:0] _4994;
    wire [64:0] _3051;
    wire [64:0] _3050;
    wire _3052;
    wire [63:0] _4993;
    wire _3049;
    wire [63:0] _4995;
    wire [63:0] _4996;
    wire _4992;
    wire [63:0] _4997;
    wire [63:0] _329;
    reg [63:0] _674;
    wire [64:0] _3066;
    wire _3068;
    wire [63:0] _4999;
    wire _3065;
    wire [63:0] _5001;
    wire [63:0] _5002;
    wire _4998;
    wire [63:0] _5003;
    wire [63:0] _330;
    reg [63:0] _671;
    wire [64:0] _3089;
    wire _3091;
    wire [63:0] _5006;
    wire [64:0] _3083;
    wire [64:0] _3082;
    wire _3084;
    wire [63:0] _5005;
    wire _3081;
    wire [63:0] _5007;
    wire [63:0] _5008;
    wire _5004;
    wire [63:0] _5009;
    wire [63:0] _331;
    reg [63:0] _668;
    wire [64:0] _3098;
    wire _3100;
    wire [63:0] _5011;
    wire _3097;
    wire [63:0] _5013;
    wire [63:0] _5014;
    wire _5010;
    wire [63:0] _5015;
    wire [63:0] _332;
    reg [63:0] _665;
    wire [64:0] _3121;
    wire _3123;
    wire [63:0] _5018;
    wire [64:0] _3115;
    wire [64:0] _3114;
    wire _3116;
    wire [63:0] _5017;
    wire _3113;
    wire [63:0] _5019;
    wire [63:0] _5020;
    wire _5016;
    wire [63:0] _5021;
    wire [63:0] _333;
    reg [63:0] _662;
    wire [64:0] _3130;
    wire _3132;
    wire [63:0] _5023;
    wire _3129;
    wire [63:0] _5025;
    wire [63:0] _5026;
    wire _5022;
    wire [63:0] _5027;
    wire [63:0] _334;
    reg [63:0] _659;
    wire [64:0] _3153;
    wire _3155;
    wire [63:0] _5030;
    wire [64:0] _3147;
    wire [64:0] _3146;
    wire _3148;
    wire [63:0] _5029;
    wire _3145;
    wire [63:0] _5031;
    wire [63:0] _5032;
    wire _5028;
    wire [63:0] _5033;
    wire [63:0] _335;
    reg [63:0] _656;
    wire [64:0] _3162;
    wire _3164;
    wire [63:0] _5035;
    wire _3161;
    wire [63:0] _5037;
    wire [63:0] _5038;
    wire _5034;
    wire [63:0] _5039;
    wire [63:0] _336;
    reg [63:0] _653;
    wire [64:0] _3185;
    wire _3187;
    wire [63:0] _5042;
    wire [64:0] _3179;
    wire [64:0] _3178;
    wire _3180;
    wire [63:0] _5041;
    wire _3177;
    wire [63:0] _5043;
    wire [63:0] _5044;
    wire _5040;
    wire [63:0] _5045;
    wire [63:0] _337;
    reg [63:0] _650;
    wire [64:0] _3194;
    wire _3196;
    wire [63:0] _5047;
    wire _3193;
    wire [63:0] _5049;
    wire [63:0] _5050;
    wire _5046;
    wire [63:0] _5051;
    wire [63:0] _338;
    reg [63:0] _647;
    wire [64:0] _3217;
    wire _3219;
    wire [63:0] _5054;
    wire [64:0] _3211;
    wire [64:0] _3210;
    wire _3212;
    wire [63:0] _5053;
    wire _3209;
    wire [63:0] _5055;
    wire [63:0] _5056;
    wire _5052;
    wire [63:0] _5057;
    wire [63:0] _339;
    reg [63:0] _644;
    wire [64:0] _3226;
    wire _3228;
    wire [63:0] _5059;
    wire _3225;
    wire [63:0] _5061;
    wire [63:0] _5062;
    wire _5058;
    wire [63:0] _5063;
    wire [63:0] _340;
    reg [63:0] _641;
    wire [64:0] _3249;
    wire _3251;
    wire [63:0] _5066;
    wire [64:0] _3243;
    wire [64:0] _3242;
    wire _3244;
    wire [63:0] _5065;
    wire _3241;
    wire [63:0] _5067;
    wire [63:0] _5068;
    wire _5064;
    wire [63:0] _5069;
    wire [63:0] _341;
    reg [63:0] _638;
    wire [64:0] _3258;
    wire _3260;
    wire [63:0] _5071;
    wire _3257;
    wire [63:0] _5073;
    wire [63:0] _5074;
    wire _5070;
    wire [63:0] _5075;
    wire [63:0] _342;
    reg [63:0] _635;
    wire [64:0] _3281;
    wire _3283;
    wire [63:0] _5078;
    wire [64:0] _3275;
    wire [64:0] _3274;
    wire _3276;
    wire [63:0] _5077;
    wire _3273;
    wire [63:0] _5079;
    wire [63:0] _5080;
    wire _5076;
    wire [63:0] _5081;
    wire [63:0] _343;
    reg [63:0] _632;
    wire [64:0] _3290;
    wire _3292;
    wire [63:0] _5083;
    wire _3289;
    wire [63:0] _5085;
    wire [63:0] _5086;
    wire _5082;
    wire [63:0] _5087;
    wire [63:0] _344;
    reg [63:0] _629;
    wire [64:0] _3313;
    wire _3315;
    wire [63:0] _5090;
    wire [64:0] _3307;
    wire [64:0] _3306;
    wire _3308;
    wire [63:0] _5089;
    wire _3305;
    wire [63:0] _5091;
    wire [63:0] _5092;
    wire _5088;
    wire [63:0] _5093;
    wire [63:0] _345;
    reg [63:0] _626;
    wire [64:0] _3322;
    wire _3324;
    wire [63:0] _5095;
    wire _3321;
    wire [63:0] _5097;
    wire [63:0] _5098;
    wire _5094;
    wire [63:0] _5099;
    wire [63:0] _346;
    reg [63:0] _623;
    wire [64:0] _3345;
    wire _3347;
    wire [63:0] _5102;
    wire [64:0] _3339;
    wire [64:0] _3338;
    wire _3340;
    wire [63:0] _5101;
    wire _3337;
    wire [63:0] _5103;
    wire [63:0] _5104;
    wire _5100;
    wire [63:0] _5105;
    wire [63:0] _347;
    reg [63:0] _620;
    wire [64:0] _3354;
    wire _3356;
    wire [63:0] _5107;
    wire _3353;
    wire [63:0] _5109;
    wire [63:0] _5110;
    wire _5106;
    wire [63:0] _5111;
    wire [63:0] _348;
    reg [63:0] _617;
    wire [64:0] _3377;
    wire _3379;
    wire [63:0] _5114;
    wire [64:0] _3371;
    wire [64:0] _3370;
    wire _3372;
    wire [63:0] _5113;
    wire _3369;
    wire [63:0] _5115;
    wire [63:0] _5116;
    wire _5112;
    wire [63:0] _5117;
    wire [63:0] _349;
    reg [63:0] _614;
    wire [64:0] _3386;
    wire _3388;
    wire [63:0] _5119;
    wire _3385;
    wire [63:0] _5121;
    wire [63:0] _5122;
    wire _5118;
    wire [63:0] _5123;
    wire [63:0] _350;
    reg [63:0] _611;
    wire [64:0] _3409;
    wire _3411;
    wire [63:0] _5126;
    wire [64:0] _3403;
    wire [64:0] _3402;
    wire _3404;
    wire [63:0] _5125;
    wire _3401;
    wire [63:0] _5127;
    wire [63:0] _5128;
    wire _5124;
    wire [63:0] _5129;
    wire [63:0] _351;
    reg [63:0] _608;
    wire [64:0] _3418;
    wire _3420;
    wire [63:0] _5131;
    wire _3417;
    wire [63:0] _5133;
    wire [63:0] _5134;
    wire _5130;
    wire [63:0] _5135;
    wire [63:0] _352;
    reg [63:0] _605;
    wire [64:0] _3441;
    wire _3443;
    wire [63:0] _5138;
    wire [64:0] _3435;
    wire [64:0] _3434;
    wire _3436;
    wire [63:0] _5137;
    wire _3433;
    wire [63:0] _5139;
    wire [63:0] _5140;
    wire _5136;
    wire [63:0] _5141;
    wire [63:0] _353;
    reg [63:0] _602;
    wire [64:0] _3450;
    wire _3452;
    wire [63:0] _5143;
    wire _3449;
    wire [63:0] _5145;
    wire [63:0] _5146;
    wire _5142;
    wire [63:0] _5147;
    wire [63:0] _354;
    reg [63:0] _599;
    wire [64:0] _3473;
    wire _3475;
    wire [63:0] _5150;
    wire [64:0] _3467;
    wire [64:0] _3466;
    wire _3468;
    wire [63:0] _5149;
    wire _3465;
    wire [63:0] _5151;
    wire [63:0] _5152;
    wire _5148;
    wire [63:0] _5153;
    wire [63:0] _355;
    reg [63:0] _596;
    wire [64:0] _3482;
    wire _3484;
    wire [63:0] _5155;
    wire _3481;
    wire [63:0] _5157;
    wire [63:0] _5158;
    wire _5154;
    wire [63:0] _5159;
    wire [63:0] _356;
    reg [63:0] _593;
    wire [64:0] _3505;
    wire _3507;
    wire [63:0] _5162;
    wire [64:0] _3499;
    wire [64:0] _3498;
    wire _3500;
    wire [63:0] _5161;
    wire _3497;
    wire [63:0] _5163;
    wire [63:0] _5164;
    wire _5160;
    wire [63:0] _5165;
    wire [63:0] _357;
    reg [63:0] _590;
    wire [64:0] _3514;
    wire _3516;
    wire [63:0] _5167;
    wire _3513;
    wire [63:0] _5169;
    wire [63:0] _5170;
    wire _5166;
    wire [63:0] _5171;
    wire [63:0] _358;
    reg [63:0] _587;
    wire [64:0] _3537;
    wire _3539;
    wire [63:0] _5174;
    wire [64:0] _3531;
    wire [64:0] _3530;
    wire _3532;
    wire [63:0] _5173;
    wire _3529;
    wire [63:0] _5175;
    wire [63:0] _5176;
    wire _5172;
    wire [63:0] _5177;
    wire [63:0] _359;
    reg [63:0] _584;
    wire [64:0] _3546;
    wire _3548;
    wire [63:0] _5179;
    wire _3545;
    wire [63:0] _5181;
    wire [63:0] _5182;
    wire _5178;
    wire [63:0] _5183;
    wire [63:0] _360;
    reg [63:0] _581;
    wire [64:0] _3569;
    wire _3571;
    wire [63:0] _5186;
    wire [64:0] _3563;
    wire [64:0] _3562;
    wire _3564;
    wire [63:0] _5185;
    wire _3561;
    wire [63:0] _5187;
    wire [63:0] _5188;
    wire _5184;
    wire [63:0] _5189;
    wire [63:0] _361;
    reg [63:0] _578;
    wire [64:0] _3578;
    wire _3580;
    wire [63:0] _5191;
    wire _3577;
    wire [63:0] _5193;
    wire [63:0] _5194;
    wire _5190;
    wire [63:0] _5195;
    wire [63:0] _362;
    reg [63:0] _575;
    wire [64:0] _3601;
    wire _3603;
    wire [63:0] _5198;
    wire [64:0] _3595;
    wire [64:0] _3594;
    wire _3596;
    wire [63:0] _5197;
    wire _3593;
    wire [63:0] _5199;
    wire [63:0] _5200;
    wire _5196;
    wire [63:0] _5201;
    wire [63:0] _363;
    reg [63:0] _572;
    wire [64:0] _3610;
    wire _3612;
    wire [63:0] _5203;
    wire _3609;
    wire [63:0] _5205;
    wire [63:0] _5206;
    wire _5202;
    wire [63:0] _5207;
    wire [63:0] _364;
    reg [63:0] _569;
    wire [64:0] _3633;
    wire _3635;
    wire [63:0] _5210;
    wire [64:0] _3627;
    wire [64:0] _3626;
    wire _3628;
    wire [63:0] _5209;
    wire _3625;
    wire [63:0] _5211;
    wire [63:0] _5212;
    wire _5208;
    wire [63:0] _5213;
    wire [63:0] _365;
    reg [63:0] _566;
    wire [64:0] _3642;
    wire _3644;
    wire [63:0] _5215;
    wire _3641;
    wire [63:0] _5217;
    wire [63:0] _5218;
    wire _5214;
    wire [63:0] _5219;
    wire [63:0] _366;
    reg [63:0] _563;
    wire [64:0] _3665;
    wire _3667;
    wire [63:0] _5222;
    wire [64:0] _3659;
    wire [64:0] _3658;
    wire _3660;
    wire [63:0] _5221;
    wire _3657;
    wire [63:0] _5223;
    wire [63:0] _5224;
    wire _5220;
    wire [63:0] _5225;
    wire [63:0] _367;
    reg [63:0] _560;
    wire [64:0] _3674;
    wire _3676;
    wire [63:0] _5227;
    wire _3673;
    wire [63:0] _5229;
    wire [63:0] _5230;
    wire _5226;
    wire [63:0] _5231;
    wire [63:0] _368;
    reg [63:0] _557;
    wire [64:0] _3697;
    wire _3699;
    wire [63:0] _5234;
    wire [64:0] _3691;
    wire [64:0] _3690;
    wire _3692;
    wire [63:0] _5233;
    wire _3689;
    wire [63:0] _5235;
    wire [63:0] _5236;
    wire _5232;
    wire [63:0] _5237;
    wire [63:0] _369;
    reg [63:0] _554;
    wire [64:0] _3706;
    wire _3708;
    wire [63:0] _5239;
    wire _3705;
    wire [63:0] _5241;
    wire [63:0] _5242;
    wire _5238;
    wire [63:0] _5243;
    wire [63:0] _370;
    reg [63:0] _551;
    wire [64:0] _3729;
    wire _3731;
    wire [63:0] _5246;
    wire [64:0] _3723;
    wire [64:0] _3722;
    wire _3724;
    wire [63:0] _5245;
    wire _3721;
    wire [63:0] _5247;
    wire [63:0] _5248;
    wire _5244;
    wire [63:0] _5249;
    wire [63:0] _371;
    reg [63:0] _548;
    wire [64:0] _3738;
    wire _3740;
    wire [63:0] _5251;
    wire _3737;
    wire [63:0] _5253;
    wire [63:0] _5254;
    wire _5250;
    wire [63:0] _5255;
    wire [63:0] _372;
    reg [63:0] _545;
    wire [64:0] _3761;
    wire _3763;
    wire [63:0] _5258;
    wire [64:0] _3755;
    wire [64:0] _3754;
    wire _3756;
    wire [63:0] _5257;
    wire _3753;
    wire [63:0] _5259;
    wire [63:0] _5260;
    wire _5256;
    wire [63:0] _5261;
    wire [63:0] _373;
    reg [63:0] _542;
    wire [64:0] _3770;
    wire _3772;
    wire [63:0] _5263;
    wire _3769;
    wire [63:0] _5265;
    wire [63:0] _5266;
    wire _5262;
    wire [63:0] _5267;
    wire [63:0] _374;
    reg [63:0] _539;
    wire [64:0] _3793;
    wire _3795;
    wire [63:0] _5270;
    wire [64:0] _3787;
    wire [64:0] _3786;
    wire _3788;
    wire [63:0] _5269;
    wire _3785;
    wire [63:0] _5271;
    wire [63:0] _5272;
    wire _5268;
    wire [63:0] _5273;
    wire [63:0] _375;
    reg [63:0] _536;
    wire [64:0] _3802;
    wire _3804;
    wire [63:0] _5275;
    wire _3801;
    wire [63:0] _5277;
    wire [63:0] _5278;
    wire _5274;
    wire [63:0] _5279;
    wire [63:0] _376;
    reg [63:0] _533;
    wire [64:0] _3825;
    wire _3827;
    wire [63:0] _5282;
    wire [64:0] _3819;
    wire [64:0] _3818;
    wire _3820;
    wire [63:0] _5281;
    wire _3817;
    wire [63:0] _5283;
    wire [63:0] _5284;
    wire _5280;
    wire [63:0] _5285;
    wire [63:0] _377;
    reg [63:0] _530;
    wire [64:0] _3834;
    wire _3836;
    wire [63:0] _5287;
    wire _3833;
    wire [63:0] _5289;
    wire [63:0] _5290;
    wire _5286;
    wire [63:0] _5291;
    wire [63:0] _378;
    reg [63:0] _527;
    wire [64:0] _3857;
    wire _3859;
    wire [63:0] _5294;
    wire [64:0] _3851;
    wire [64:0] _3850;
    wire _3852;
    wire [63:0] _5293;
    wire _3849;
    wire [63:0] _5295;
    wire [63:0] _5296;
    wire _5292;
    wire [63:0] _5297;
    wire [63:0] _379;
    reg [63:0] _524;
    wire [64:0] _3866;
    wire _3868;
    wire [63:0] _5299;
    wire _3865;
    wire [63:0] _5301;
    wire [63:0] _5302;
    wire _5298;
    wire [63:0] _5303;
    wire [63:0] _380;
    reg [63:0] _521;
    wire [64:0] _3889;
    wire _3891;
    wire [63:0] _5306;
    wire [64:0] _3883;
    wire [64:0] _3882;
    wire _3884;
    wire [63:0] _5305;
    wire _3881;
    wire [63:0] _5307;
    wire [63:0] _5308;
    wire _5304;
    wire [63:0] _5309;
    wire [63:0] _381;
    reg [63:0] _518;
    wire [64:0] _3898;
    wire _3900;
    wire [63:0] _5311;
    wire _3897;
    wire [63:0] _5313;
    wire [63:0] _5314;
    wire _5310;
    wire [63:0] _5315;
    wire [63:0] _382;
    reg [63:0] _515;
    wire [64:0] _3921;
    wire _3923;
    wire [63:0] _5318;
    wire [64:0] _3915;
    wire [64:0] _3914;
    wire _3916;
    wire [63:0] _5317;
    wire _3913;
    wire [63:0] _5319;
    wire [63:0] _5320;
    wire _5316;
    wire [63:0] _5321;
    wire [63:0] _383;
    reg [63:0] _512;
    wire [64:0] _3930;
    wire _3932;
    wire [63:0] _5323;
    wire _3929;
    wire [63:0] _5325;
    wire [63:0] _5326;
    wire _5322;
    wire [63:0] _5327;
    wire [63:0] _384;
    reg [63:0] _509;
    wire [64:0] _3953;
    wire _3955;
    wire [63:0] _5330;
    wire [64:0] _3947;
    wire [64:0] _3946;
    wire _3948;
    wire [63:0] _5329;
    wire _3945;
    wire [63:0] _5331;
    wire [63:0] _5332;
    wire _5328;
    wire [63:0] _5333;
    wire [63:0] _385;
    reg [63:0] _506;
    wire [64:0] _3962;
    wire _3964;
    wire [63:0] _5335;
    wire _3961;
    wire [63:0] _5337;
    wire [63:0] _5338;
    wire _5334;
    wire [63:0] _5339;
    wire [63:0] _386;
    reg [63:0] _503;
    wire [64:0] _3985;
    wire _3987;
    wire [63:0] _5342;
    wire [64:0] _3979;
    wire [64:0] _3978;
    wire _3980;
    wire [63:0] _5341;
    wire _3977;
    wire [63:0] _5343;
    wire [63:0] _5344;
    wire _5340;
    wire [63:0] _5345;
    wire [63:0] _387;
    reg [63:0] _500;
    wire [64:0] _3994;
    wire _3996;
    wire [63:0] _5347;
    wire _3993;
    wire [63:0] _5349;
    wire [63:0] _5350;
    wire _5346;
    wire [63:0] _5351;
    wire [63:0] _388;
    reg [63:0] _497;
    wire [64:0] _4017;
    wire _4019;
    wire [63:0] _5354;
    wire [64:0] _4011;
    wire [64:0] _4010;
    wire _4012;
    wire [63:0] _5353;
    wire _4009;
    wire [63:0] _5355;
    wire [63:0] _5356;
    wire _5352;
    wire [63:0] _5357;
    wire [63:0] _389;
    reg [63:0] _494;
    wire [64:0] _4026;
    wire _4028;
    wire [63:0] _5359;
    wire _4025;
    wire [63:0] _5361;
    wire [63:0] _5362;
    wire _5358;
    wire [63:0] _5363;
    wire [63:0] _390;
    reg [63:0] _491;
    wire [64:0] _4049;
    wire _4051;
    wire [63:0] _5366;
    wire [64:0] _4043;
    wire [64:0] _4042;
    wire _4044;
    wire [63:0] _5365;
    wire _4041;
    wire [63:0] _5367;
    wire [63:0] _5368;
    wire _5364;
    wire [63:0] _5369;
    wire [63:0] _391;
    reg [63:0] _488;
    wire [64:0] _4058;
    wire _4060;
    wire [63:0] _5371;
    wire _4057;
    wire [63:0] _5373;
    wire [63:0] _5374;
    wire _5370;
    wire [63:0] _5375;
    wire [63:0] _392;
    reg [63:0] _485;
    wire [64:0] _4081;
    wire _4083;
    wire [63:0] _5378;
    wire [64:0] _4075;
    wire [64:0] _4074;
    wire _4076;
    wire [63:0] _5377;
    wire _4073;
    wire [63:0] _5379;
    wire [63:0] _5380;
    wire _5376;
    wire [63:0] _5381;
    wire [63:0] _393;
    reg [63:0] _482;
    wire [64:0] _4090;
    wire _4092;
    wire [63:0] _5383;
    wire _4089;
    wire [63:0] _5385;
    wire [63:0] _5386;
    wire _5382;
    wire [63:0] _5387;
    wire [63:0] _394;
    reg [63:0] _479;
    wire [64:0] _4113;
    wire _4115;
    wire [63:0] _5390;
    wire [64:0] _4107;
    wire [64:0] _4106;
    wire _4108;
    wire [63:0] _5389;
    wire _4105;
    wire [63:0] _5391;
    wire [63:0] _5392;
    wire _5388;
    wire [63:0] _5393;
    wire [63:0] _395;
    reg [63:0] _476;
    wire [64:0] _4122;
    wire _4124;
    wire [63:0] _5395;
    wire _4121;
    wire [63:0] _5397;
    wire [63:0] _5398;
    wire _5394;
    wire [63:0] _5399;
    wire [63:0] _396;
    reg [63:0] _473;
    wire [64:0] _4145;
    wire _4147;
    wire [63:0] _5402;
    wire [64:0] _4139;
    wire [64:0] _4138;
    wire _4140;
    wire [63:0] _5401;
    wire _4137;
    wire [63:0] _5403;
    wire [63:0] _5404;
    wire _5400;
    wire [63:0] _5405;
    wire [63:0] _397;
    reg [63:0] _470;
    wire [64:0] _4154;
    wire _4156;
    wire [63:0] _5407;
    wire _4153;
    wire [63:0] _5409;
    wire [63:0] _5410;
    wire _5406;
    wire [63:0] _5411;
    wire [63:0] _398;
    reg [63:0] _467;
    wire [64:0] _4177;
    wire _4179;
    wire [63:0] _5414;
    wire [64:0] _4171;
    wire [64:0] _4170;
    wire _4172;
    wire [63:0] _5413;
    wire _4169;
    wire [63:0] _5415;
    wire [63:0] _5416;
    wire _5412;
    wire [63:0] _5417;
    wire [63:0] _399;
    reg [63:0] _464;
    wire [64:0] _4186;
    wire _4188;
    wire [63:0] _5419;
    wire _4185;
    wire [63:0] _5421;
    wire [63:0] _5422;
    wire _5418;
    wire [63:0] _5423;
    wire [63:0] _400;
    reg [63:0] _461;
    wire [64:0] _4209;
    wire _4211;
    wire [63:0] _5426;
    wire [64:0] _4203;
    wire [64:0] _4202;
    wire _4204;
    wire [63:0] _5425;
    wire _4201;
    wire [63:0] _5427;
    wire [63:0] _5428;
    wire _5424;
    wire [63:0] _5429;
    wire [63:0] _401;
    reg [63:0] _458;
    wire [64:0] _4218;
    wire _4220;
    wire [63:0] _5431;
    wire _4217;
    wire [63:0] _5433;
    wire [63:0] _5434;
    wire _5430;
    wire [63:0] _5435;
    wire [63:0] _402;
    reg [63:0] _455;
    wire [64:0] _4241;
    wire _4243;
    wire [63:0] _5451;
    wire [63:0] _404;
    wire [64:0] _5443;
    wire [64:0] _5442;
    wire _5444;
    wire [63:0] _5445;
    wire [63:0] _5441;
    wire [63:0] _5446;
    wire [63:0] _5447;
    wire _5436;
    wire [63:0] _5448;
    wire [63:0] _405;
    reg [63:0] _449;
    wire [64:0] _4235;
    wire [64:0] _4234;
    wire _4236;
    wire [63:0] _5450;
    wire _4233;
    wire [63:0] _5452;
    wire [63:0] _5453;
    wire _5449;
    wire [63:0] _5454;
    wire [63:0] _406;
    reg [63:0] _452;
    wire [64:0] _5438;
    wire _5440;
    wire [63:0] _5456;
    wire _5437;
    wire [63:0] _5458;
    wire [63:0] _5459;
    wire _408;
    wire _1055;
    wire _5455;
    wire [63:0] _5460;
    wire [63:0] _409;
    reg [63:0] _4239;
    reg [63:0] _5462;
    wire _5461;
    wire [63:0] _5467;
    wire [63:0] _5468;
    wire [63:0] _410;
    reg [63:0] _440;
    wire [63:0] _442;
    wire [64:0] _443;
    wire _1049;
    wire _1050;
    wire _5488;
    wire _5489;
    wire _435;
    wire _5473;
    wire _5474;
    wire _411;
    reg _436;
    wire vdd;
    wire [1:0] _424;
    wire [1:0] _427;
    wire [16:0] _5470;
    wire [15:0] _445;
    wire [15:0] _5475;
    wire [15:0] _5476;
    wire [15:0] _412;
    reg [15:0] _446;
    wire [16:0] _5469;
    wire _5471;
    wire _5472;
    wire [1:0] _5485;
    wire [1:0] _429;
    wire _1058;
    wire _414;
    wire _416;
    wire [15:0] _5478;
    wire [15:0] _417;
    reg [15:0] _1064;
    wire gnd;
    wire [16:0] _5480;
    wire _5482;
    wire _5483;
    wire [1:0] _5484;
    wire [1:0] _1057;
    wire _419;
    wire [1:0] _5479;
    reg [1:0] _5486;
    wire [1:0] _420;
    reg [1:0] _426;
    wire _430;
    wire _5487;
    wire _5490;
    wire [63:0] _5498;
    wire [63:0] _421;
    reg [63:0] _5493;
    assign _428 = _426 == _427;
    assign _5492 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _5495 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    assign _1051 = _436 & _1050;
    assign _1052 = _1051 ? _433 : _1047;
    assign _1053 = _430 ? _1052 : _433;
    assign _3 = _1053;
    always @(posedge _416) begin
        if (_414)
            _433 <= _5492;
        else
            _433 <= _3;
    end
    assign _5494 = _440 - _433;
    assign _5496 = _5494 + _5495;
    assign _5497 = _5493 + _5496;
    always @* begin
        case (_446)
        0:
            _1047 <= _449;
        1:
            _1047 <= _452;
        2:
            _1047 <= _455;
        3:
            _1047 <= _458;
        4:
            _1047 <= _461;
        5:
            _1047 <= _464;
        6:
            _1047 <= _467;
        7:
            _1047 <= _470;
        8:
            _1047 <= _473;
        9:
            _1047 <= _476;
        10:
            _1047 <= _479;
        11:
            _1047 <= _482;
        12:
            _1047 <= _485;
        13:
            _1047 <= _488;
        14:
            _1047 <= _491;
        15:
            _1047 <= _494;
        16:
            _1047 <= _497;
        17:
            _1047 <= _500;
        18:
            _1047 <= _503;
        19:
            _1047 <= _506;
        20:
            _1047 <= _509;
        21:
            _1047 <= _512;
        22:
            _1047 <= _515;
        23:
            _1047 <= _518;
        24:
            _1047 <= _521;
        25:
            _1047 <= _524;
        26:
            _1047 <= _527;
        27:
            _1047 <= _530;
        28:
            _1047 <= _533;
        29:
            _1047 <= _536;
        30:
            _1047 <= _539;
        31:
            _1047 <= _542;
        32:
            _1047 <= _545;
        33:
            _1047 <= _548;
        34:
            _1047 <= _551;
        35:
            _1047 <= _554;
        36:
            _1047 <= _557;
        37:
            _1047 <= _560;
        38:
            _1047 <= _563;
        39:
            _1047 <= _566;
        40:
            _1047 <= _569;
        41:
            _1047 <= _572;
        42:
            _1047 <= _575;
        43:
            _1047 <= _578;
        44:
            _1047 <= _581;
        45:
            _1047 <= _584;
        46:
            _1047 <= _587;
        47:
            _1047 <= _590;
        48:
            _1047 <= _593;
        49:
            _1047 <= _596;
        50:
            _1047 <= _599;
        51:
            _1047 <= _602;
        52:
            _1047 <= _605;
        53:
            _1047 <= _608;
        54:
            _1047 <= _611;
        55:
            _1047 <= _614;
        56:
            _1047 <= _617;
        57:
            _1047 <= _620;
        58:
            _1047 <= _623;
        59:
            _1047 <= _626;
        60:
            _1047 <= _629;
        61:
            _1047 <= _632;
        62:
            _1047 <= _635;
        63:
            _1047 <= _638;
        64:
            _1047 <= _641;
        65:
            _1047 <= _644;
        66:
            _1047 <= _647;
        67:
            _1047 <= _650;
        68:
            _1047 <= _653;
        69:
            _1047 <= _656;
        70:
            _1047 <= _659;
        71:
            _1047 <= _662;
        72:
            _1047 <= _665;
        73:
            _1047 <= _668;
        74:
            _1047 <= _671;
        75:
            _1047 <= _674;
        76:
            _1047 <= _677;
        77:
            _1047 <= _680;
        78:
            _1047 <= _683;
        79:
            _1047 <= _686;
        80:
            _1047 <= _689;
        81:
            _1047 <= _692;
        82:
            _1047 <= _695;
        83:
            _1047 <= _698;
        84:
            _1047 <= _701;
        85:
            _1047 <= _704;
        86:
            _1047 <= _707;
        87:
            _1047 <= _710;
        88:
            _1047 <= _713;
        89:
            _1047 <= _716;
        90:
            _1047 <= _719;
        91:
            _1047 <= _722;
        92:
            _1047 <= _725;
        93:
            _1047 <= _728;
        94:
            _1047 <= _731;
        95:
            _1047 <= _734;
        96:
            _1047 <= _737;
        97:
            _1047 <= _740;
        98:
            _1047 <= _743;
        99:
            _1047 <= _746;
        100:
            _1047 <= _749;
        101:
            _1047 <= _752;
        102:
            _1047 <= _755;
        103:
            _1047 <= _758;
        104:
            _1047 <= _761;
        105:
            _1047 <= _764;
        106:
            _1047 <= _767;
        107:
            _1047 <= _770;
        108:
            _1047 <= _773;
        109:
            _1047 <= _776;
        110:
            _1047 <= _779;
        111:
            _1047 <= _782;
        112:
            _1047 <= _785;
        113:
            _1047 <= _788;
        114:
            _1047 <= _791;
        115:
            _1047 <= _794;
        116:
            _1047 <= _797;
        117:
            _1047 <= _800;
        118:
            _1047 <= _803;
        119:
            _1047 <= _806;
        120:
            _1047 <= _809;
        121:
            _1047 <= _812;
        122:
            _1047 <= _815;
        123:
            _1047 <= _818;
        124:
            _1047 <= _821;
        125:
            _1047 <= _824;
        126:
            _1047 <= _827;
        127:
            _1047 <= _830;
        128:
            _1047 <= _833;
        129:
            _1047 <= _836;
        130:
            _1047 <= _839;
        131:
            _1047 <= _842;
        132:
            _1047 <= _845;
        133:
            _1047 <= _848;
        134:
            _1047 <= _851;
        135:
            _1047 <= _854;
        136:
            _1047 <= _857;
        137:
            _1047 <= _860;
        138:
            _1047 <= _863;
        139:
            _1047 <= _866;
        140:
            _1047 <= _869;
        141:
            _1047 <= _872;
        142:
            _1047 <= _875;
        143:
            _1047 <= _878;
        144:
            _1047 <= _881;
        145:
            _1047 <= _884;
        146:
            _1047 <= _887;
        147:
            _1047 <= _890;
        148:
            _1047 <= _893;
        149:
            _1047 <= _896;
        150:
            _1047 <= _899;
        151:
            _1047 <= _902;
        152:
            _1047 <= _905;
        153:
            _1047 <= _908;
        154:
            _1047 <= _911;
        155:
            _1047 <= _914;
        156:
            _1047 <= _917;
        157:
            _1047 <= _920;
        158:
            _1047 <= _923;
        159:
            _1047 <= _926;
        160:
            _1047 <= _929;
        161:
            _1047 <= _932;
        162:
            _1047 <= _935;
        163:
            _1047 <= _938;
        164:
            _1047 <= _941;
        165:
            _1047 <= _944;
        166:
            _1047 <= _947;
        167:
            _1047 <= _950;
        168:
            _1047 <= _953;
        169:
            _1047 <= _956;
        170:
            _1047 <= _959;
        171:
            _1047 <= _962;
        172:
            _1047 <= _965;
        173:
            _1047 <= _968;
        174:
            _1047 <= _971;
        175:
            _1047 <= _974;
        176:
            _1047 <= _977;
        177:
            _1047 <= _980;
        178:
            _1047 <= _983;
        179:
            _1047 <= _986;
        180:
            _1047 <= _989;
        181:
            _1047 <= _992;
        182:
            _1047 <= _995;
        183:
            _1047 <= _998;
        184:
            _1047 <= _1001;
        185:
            _1047 <= _1004;
        186:
            _1047 <= _1007;
        187:
            _1047 <= _1010;
        188:
            _1047 <= _1013;
        189:
            _1047 <= _1016;
        190:
            _1047 <= _1019;
        191:
            _1047 <= _1022;
        192:
            _1047 <= _1025;
        193:
            _1047 <= _1028;
        194:
            _1047 <= _1031;
        195:
            _1047 <= _1034;
        196:
            _1047 <= _1037;
        197:
            _1047 <= _1040;
        198:
            _1047 <= _1043;
        default:
            _1047 <= _1046;
        endcase
    end
    assign _1048 = { gnd,
                     _1047 };
    assign _5464 = { gnd,
                     _5462 };
    assign _5463 = { gnd,
                     _440 };
    assign _5465 = _5463 < _5464;
    assign _5466 = _5465 ? _5462 : _440;
    assign _5 = wr_end;
    assign _5457 = _5444 ? _4239 : _4239;
    assign _4228 = _4224 ? _4227 : _4207;
    assign _4196 = _4192 ? _4195 : _4175;
    assign _4164 = _4160 ? _4163 : _4143;
    assign _4132 = _4128 ? _4131 : _4111;
    assign _4100 = _4096 ? _4099 : _4079;
    assign _4068 = _4064 ? _4067 : _4047;
    assign _4036 = _4032 ? _4035 : _4015;
    assign _4004 = _4000 ? _4003 : _3983;
    assign _3972 = _3968 ? _3971 : _3951;
    assign _3940 = _3936 ? _3939 : _3919;
    assign _3908 = _3904 ? _3907 : _3887;
    assign _3876 = _3872 ? _3875 : _3855;
    assign _3844 = _3840 ? _3843 : _3823;
    assign _3812 = _3808 ? _3811 : _3791;
    assign _3780 = _3776 ? _3779 : _3759;
    assign _3748 = _3744 ? _3747 : _3727;
    assign _3716 = _3712 ? _3715 : _3695;
    assign _3684 = _3680 ? _3683 : _3663;
    assign _3652 = _3648 ? _3651 : _3631;
    assign _3620 = _3616 ? _3619 : _3599;
    assign _3588 = _3584 ? _3587 : _3567;
    assign _3556 = _3552 ? _3555 : _3535;
    assign _3524 = _3520 ? _3523 : _3503;
    assign _3492 = _3488 ? _3491 : _3471;
    assign _3460 = _3456 ? _3459 : _3439;
    assign _3428 = _3424 ? _3427 : _3407;
    assign _3396 = _3392 ? _3395 : _3375;
    assign _3364 = _3360 ? _3363 : _3343;
    assign _3332 = _3328 ? _3331 : _3311;
    assign _3300 = _3296 ? _3299 : _3279;
    assign _3268 = _3264 ? _3267 : _3247;
    assign _3236 = _3232 ? _3235 : _3215;
    assign _3204 = _3200 ? _3203 : _3183;
    assign _3172 = _3168 ? _3171 : _3151;
    assign _3140 = _3136 ? _3139 : _3119;
    assign _3108 = _3104 ? _3107 : _3087;
    assign _3076 = _3072 ? _3075 : _3055;
    assign _3044 = _3040 ? _3043 : _3023;
    assign _3012 = _3008 ? _3011 : _2991;
    assign _2980 = _2976 ? _2979 : _2959;
    assign _2948 = _2944 ? _2947 : _2927;
    assign _2916 = _2912 ? _2915 : _2895;
    assign _2884 = _2880 ? _2883 : _2863;
    assign _2852 = _2848 ? _2851 : _2831;
    assign _2820 = _2816 ? _2819 : _2799;
    assign _2788 = _2784 ? _2787 : _2767;
    assign _2756 = _2752 ? _2755 : _2735;
    assign _2724 = _2720 ? _2723 : _2703;
    assign _2692 = _2688 ? _2691 : _2671;
    assign _2660 = _2656 ? _2659 : _2639;
    assign _2628 = _2624 ? _2627 : _2607;
    assign _2596 = _2592 ? _2595 : _2575;
    assign _2564 = _2560 ? _2563 : _2543;
    assign _2532 = _2528 ? _2531 : _2511;
    assign _2500 = _2496 ? _2499 : _2479;
    assign _2468 = _2464 ? _2467 : _2447;
    assign _2436 = _2432 ? _2435 : _2415;
    assign _2404 = _2400 ? _2403 : _2383;
    assign _2372 = _2368 ? _2371 : _2351;
    assign _2340 = _2336 ? _2339 : _2319;
    assign _2308 = _2304 ? _2307 : _2287;
    assign _2276 = _2272 ? _2275 : _2255;
    assign _2244 = _2240 ? _2243 : _2223;
    assign _2212 = _2208 ? _2211 : _2191;
    assign _2180 = _2176 ? _2179 : _2159;
    assign _2148 = _2144 ? _2147 : _2127;
    assign _2116 = _2112 ? _2115 : _2095;
    assign _2084 = _2080 ? _2083 : _2063;
    assign _2052 = _2048 ? _2051 : _2031;
    assign _2020 = _2016 ? _2019 : _1999;
    assign _1988 = _1984 ? _1987 : _1967;
    assign _1956 = _1952 ? _1955 : _1935;
    assign _1924 = _1920 ? _1923 : _1903;
    assign _1892 = _1888 ? _1891 : _1871;
    assign _1860 = _1856 ? _1859 : _1839;
    assign _1828 = _1824 ? _1827 : _1807;
    assign _1796 = _1792 ? _1795 : _1775;
    assign _1764 = _1760 ? _1763 : _1743;
    assign _1732 = _1728 ? _1731 : _1711;
    assign _1700 = _1696 ? _1699 : _1679;
    assign _1668 = _1664 ? _1667 : _1647;
    assign _1636 = _1632 ? _1635 : _1615;
    assign _1604 = _1600 ? _1603 : _1583;
    assign _1572 = _1568 ? _1571 : _1551;
    assign _1540 = _1536 ? _1539 : _1519;
    assign _1508 = _1504 ? _1507 : _1487;
    assign _1476 = _1472 ? _1475 : _1455;
    assign _1444 = _1440 ? _1443 : _1423;
    assign _1412 = _1408 ? _1411 : _1391;
    assign _1380 = _1376 ? _1379 : _1359;
    assign _1348 = _1344 ? _1347 : _1327;
    assign _1316 = _1312 ? _1315 : _1295;
    assign _1284 = _1280 ? _1283 : _1263;
    assign _1252 = _1248 ? _1251 : _1231;
    assign _1220 = _1216 ? _1219 : _1199;
    assign _1188 = _1184 ? _1187 : _1167;
    assign _1156 = _1152 ? _1155 : _1135;
    assign _1124 = _1120 ? _1123 : _1103;
    assign _1092 = _1088 ? _1091 : _1071;
    assign _1076 = _1075 ? _1061 : _1061;
    assign _1072 = _1068 ? _1071 : _1061;
    assign _1077 = _1065 ? _1076 : _1072;
    assign _1078 = _1058 ? _1077 : _1061;
    assign _1056 = _1055 & _408;
    assign _1079 = _1056 ? _1071 : _1078;
    assign _6 = _1079;
    always @(posedge _416) begin
        if (_414)
            _1061 <= _5492;
        else
            _1061 <= _6;
    end
    assign _1085 = _1084 ? _1061 : _1071;
    assign _1093 = _1081 ? _1092 : _1085;
    assign _1094 = _1058 ? _1093 : _1071;
    assign _1080 = _1055 & _408;
    assign _1095 = _1080 ? _1091 : _1094;
    assign _7 = _1095;
    always @(posedge _416) begin
        if (_414)
            _1071 <= _5492;
        else
            _1071 <= _7;
    end
    assign _1108 = _1107 ? _1071 : _1091;
    assign _1104 = _1100 ? _1103 : _1091;
    assign _1109 = _1097 ? _1108 : _1104;
    assign _1110 = _1058 ? _1109 : _1091;
    assign _1096 = _1055 & _408;
    assign _1111 = _1096 ? _1103 : _1110;
    assign _8 = _1111;
    always @(posedge _416) begin
        if (_414)
            _1091 <= _5492;
        else
            _1091 <= _8;
    end
    assign _1117 = _1116 ? _1091 : _1103;
    assign _1125 = _1113 ? _1124 : _1117;
    assign _1126 = _1058 ? _1125 : _1103;
    assign _1112 = _1055 & _408;
    assign _1127 = _1112 ? _1123 : _1126;
    assign _9 = _1127;
    always @(posedge _416) begin
        if (_414)
            _1103 <= _5492;
        else
            _1103 <= _9;
    end
    assign _1140 = _1139 ? _1103 : _1123;
    assign _1136 = _1132 ? _1135 : _1123;
    assign _1141 = _1129 ? _1140 : _1136;
    assign _1142 = _1058 ? _1141 : _1123;
    assign _1128 = _1055 & _408;
    assign _1143 = _1128 ? _1135 : _1142;
    assign _10 = _1143;
    always @(posedge _416) begin
        if (_414)
            _1123 <= _5492;
        else
            _1123 <= _10;
    end
    assign _1149 = _1148 ? _1123 : _1135;
    assign _1157 = _1145 ? _1156 : _1149;
    assign _1158 = _1058 ? _1157 : _1135;
    assign _1144 = _1055 & _408;
    assign _1159 = _1144 ? _1155 : _1158;
    assign _11 = _1159;
    always @(posedge _416) begin
        if (_414)
            _1135 <= _5492;
        else
            _1135 <= _11;
    end
    assign _1172 = _1171 ? _1135 : _1155;
    assign _1168 = _1164 ? _1167 : _1155;
    assign _1173 = _1161 ? _1172 : _1168;
    assign _1174 = _1058 ? _1173 : _1155;
    assign _1160 = _1055 & _408;
    assign _1175 = _1160 ? _1167 : _1174;
    assign _12 = _1175;
    always @(posedge _416) begin
        if (_414)
            _1155 <= _5492;
        else
            _1155 <= _12;
    end
    assign _1181 = _1180 ? _1155 : _1167;
    assign _1189 = _1177 ? _1188 : _1181;
    assign _1190 = _1058 ? _1189 : _1167;
    assign _1176 = _1055 & _408;
    assign _1191 = _1176 ? _1187 : _1190;
    assign _13 = _1191;
    always @(posedge _416) begin
        if (_414)
            _1167 <= _5492;
        else
            _1167 <= _13;
    end
    assign _1204 = _1203 ? _1167 : _1187;
    assign _1200 = _1196 ? _1199 : _1187;
    assign _1205 = _1193 ? _1204 : _1200;
    assign _1206 = _1058 ? _1205 : _1187;
    assign _1192 = _1055 & _408;
    assign _1207 = _1192 ? _1199 : _1206;
    assign _14 = _1207;
    always @(posedge _416) begin
        if (_414)
            _1187 <= _5492;
        else
            _1187 <= _14;
    end
    assign _1213 = _1212 ? _1187 : _1199;
    assign _1221 = _1209 ? _1220 : _1213;
    assign _1222 = _1058 ? _1221 : _1199;
    assign _1208 = _1055 & _408;
    assign _1223 = _1208 ? _1219 : _1222;
    assign _15 = _1223;
    always @(posedge _416) begin
        if (_414)
            _1199 <= _5492;
        else
            _1199 <= _15;
    end
    assign _1236 = _1235 ? _1199 : _1219;
    assign _1232 = _1228 ? _1231 : _1219;
    assign _1237 = _1225 ? _1236 : _1232;
    assign _1238 = _1058 ? _1237 : _1219;
    assign _1224 = _1055 & _408;
    assign _1239 = _1224 ? _1231 : _1238;
    assign _16 = _1239;
    always @(posedge _416) begin
        if (_414)
            _1219 <= _5492;
        else
            _1219 <= _16;
    end
    assign _1245 = _1244 ? _1219 : _1231;
    assign _1253 = _1241 ? _1252 : _1245;
    assign _1254 = _1058 ? _1253 : _1231;
    assign _1240 = _1055 & _408;
    assign _1255 = _1240 ? _1251 : _1254;
    assign _17 = _1255;
    always @(posedge _416) begin
        if (_414)
            _1231 <= _5492;
        else
            _1231 <= _17;
    end
    assign _1268 = _1267 ? _1231 : _1251;
    assign _1264 = _1260 ? _1263 : _1251;
    assign _1269 = _1257 ? _1268 : _1264;
    assign _1270 = _1058 ? _1269 : _1251;
    assign _1256 = _1055 & _408;
    assign _1271 = _1256 ? _1263 : _1270;
    assign _18 = _1271;
    always @(posedge _416) begin
        if (_414)
            _1251 <= _5492;
        else
            _1251 <= _18;
    end
    assign _1277 = _1276 ? _1251 : _1263;
    assign _1285 = _1273 ? _1284 : _1277;
    assign _1286 = _1058 ? _1285 : _1263;
    assign _1272 = _1055 & _408;
    assign _1287 = _1272 ? _1283 : _1286;
    assign _19 = _1287;
    always @(posedge _416) begin
        if (_414)
            _1263 <= _5492;
        else
            _1263 <= _19;
    end
    assign _1300 = _1299 ? _1263 : _1283;
    assign _1296 = _1292 ? _1295 : _1283;
    assign _1301 = _1289 ? _1300 : _1296;
    assign _1302 = _1058 ? _1301 : _1283;
    assign _1288 = _1055 & _408;
    assign _1303 = _1288 ? _1295 : _1302;
    assign _20 = _1303;
    always @(posedge _416) begin
        if (_414)
            _1283 <= _5492;
        else
            _1283 <= _20;
    end
    assign _1309 = _1308 ? _1283 : _1295;
    assign _1317 = _1305 ? _1316 : _1309;
    assign _1318 = _1058 ? _1317 : _1295;
    assign _1304 = _1055 & _408;
    assign _1319 = _1304 ? _1315 : _1318;
    assign _21 = _1319;
    always @(posedge _416) begin
        if (_414)
            _1295 <= _5492;
        else
            _1295 <= _21;
    end
    assign _1332 = _1331 ? _1295 : _1315;
    assign _1328 = _1324 ? _1327 : _1315;
    assign _1333 = _1321 ? _1332 : _1328;
    assign _1334 = _1058 ? _1333 : _1315;
    assign _1320 = _1055 & _408;
    assign _1335 = _1320 ? _1327 : _1334;
    assign _22 = _1335;
    always @(posedge _416) begin
        if (_414)
            _1315 <= _5492;
        else
            _1315 <= _22;
    end
    assign _1341 = _1340 ? _1315 : _1327;
    assign _1349 = _1337 ? _1348 : _1341;
    assign _1350 = _1058 ? _1349 : _1327;
    assign _1336 = _1055 & _408;
    assign _1351 = _1336 ? _1347 : _1350;
    assign _23 = _1351;
    always @(posedge _416) begin
        if (_414)
            _1327 <= _5492;
        else
            _1327 <= _23;
    end
    assign _1364 = _1363 ? _1327 : _1347;
    assign _1360 = _1356 ? _1359 : _1347;
    assign _1365 = _1353 ? _1364 : _1360;
    assign _1366 = _1058 ? _1365 : _1347;
    assign _1352 = _1055 & _408;
    assign _1367 = _1352 ? _1359 : _1366;
    assign _24 = _1367;
    always @(posedge _416) begin
        if (_414)
            _1347 <= _5492;
        else
            _1347 <= _24;
    end
    assign _1373 = _1372 ? _1347 : _1359;
    assign _1381 = _1369 ? _1380 : _1373;
    assign _1382 = _1058 ? _1381 : _1359;
    assign _1368 = _1055 & _408;
    assign _1383 = _1368 ? _1379 : _1382;
    assign _25 = _1383;
    always @(posedge _416) begin
        if (_414)
            _1359 <= _5492;
        else
            _1359 <= _25;
    end
    assign _1396 = _1395 ? _1359 : _1379;
    assign _1392 = _1388 ? _1391 : _1379;
    assign _1397 = _1385 ? _1396 : _1392;
    assign _1398 = _1058 ? _1397 : _1379;
    assign _1384 = _1055 & _408;
    assign _1399 = _1384 ? _1391 : _1398;
    assign _26 = _1399;
    always @(posedge _416) begin
        if (_414)
            _1379 <= _5492;
        else
            _1379 <= _26;
    end
    assign _1405 = _1404 ? _1379 : _1391;
    assign _1413 = _1401 ? _1412 : _1405;
    assign _1414 = _1058 ? _1413 : _1391;
    assign _1400 = _1055 & _408;
    assign _1415 = _1400 ? _1411 : _1414;
    assign _27 = _1415;
    always @(posedge _416) begin
        if (_414)
            _1391 <= _5492;
        else
            _1391 <= _27;
    end
    assign _1428 = _1427 ? _1391 : _1411;
    assign _1424 = _1420 ? _1423 : _1411;
    assign _1429 = _1417 ? _1428 : _1424;
    assign _1430 = _1058 ? _1429 : _1411;
    assign _1416 = _1055 & _408;
    assign _1431 = _1416 ? _1423 : _1430;
    assign _28 = _1431;
    always @(posedge _416) begin
        if (_414)
            _1411 <= _5492;
        else
            _1411 <= _28;
    end
    assign _1437 = _1436 ? _1411 : _1423;
    assign _1445 = _1433 ? _1444 : _1437;
    assign _1446 = _1058 ? _1445 : _1423;
    assign _1432 = _1055 & _408;
    assign _1447 = _1432 ? _1443 : _1446;
    assign _29 = _1447;
    always @(posedge _416) begin
        if (_414)
            _1423 <= _5492;
        else
            _1423 <= _29;
    end
    assign _1460 = _1459 ? _1423 : _1443;
    assign _1456 = _1452 ? _1455 : _1443;
    assign _1461 = _1449 ? _1460 : _1456;
    assign _1462 = _1058 ? _1461 : _1443;
    assign _1448 = _1055 & _408;
    assign _1463 = _1448 ? _1455 : _1462;
    assign _30 = _1463;
    always @(posedge _416) begin
        if (_414)
            _1443 <= _5492;
        else
            _1443 <= _30;
    end
    assign _1469 = _1468 ? _1443 : _1455;
    assign _1477 = _1465 ? _1476 : _1469;
    assign _1478 = _1058 ? _1477 : _1455;
    assign _1464 = _1055 & _408;
    assign _1479 = _1464 ? _1475 : _1478;
    assign _31 = _1479;
    always @(posedge _416) begin
        if (_414)
            _1455 <= _5492;
        else
            _1455 <= _31;
    end
    assign _1492 = _1491 ? _1455 : _1475;
    assign _1488 = _1484 ? _1487 : _1475;
    assign _1493 = _1481 ? _1492 : _1488;
    assign _1494 = _1058 ? _1493 : _1475;
    assign _1480 = _1055 & _408;
    assign _1495 = _1480 ? _1487 : _1494;
    assign _32 = _1495;
    always @(posedge _416) begin
        if (_414)
            _1475 <= _5492;
        else
            _1475 <= _32;
    end
    assign _1501 = _1500 ? _1475 : _1487;
    assign _1509 = _1497 ? _1508 : _1501;
    assign _1510 = _1058 ? _1509 : _1487;
    assign _1496 = _1055 & _408;
    assign _1511 = _1496 ? _1507 : _1510;
    assign _33 = _1511;
    always @(posedge _416) begin
        if (_414)
            _1487 <= _5492;
        else
            _1487 <= _33;
    end
    assign _1524 = _1523 ? _1487 : _1507;
    assign _1520 = _1516 ? _1519 : _1507;
    assign _1525 = _1513 ? _1524 : _1520;
    assign _1526 = _1058 ? _1525 : _1507;
    assign _1512 = _1055 & _408;
    assign _1527 = _1512 ? _1519 : _1526;
    assign _34 = _1527;
    always @(posedge _416) begin
        if (_414)
            _1507 <= _5492;
        else
            _1507 <= _34;
    end
    assign _1533 = _1532 ? _1507 : _1519;
    assign _1541 = _1529 ? _1540 : _1533;
    assign _1542 = _1058 ? _1541 : _1519;
    assign _1528 = _1055 & _408;
    assign _1543 = _1528 ? _1539 : _1542;
    assign _35 = _1543;
    always @(posedge _416) begin
        if (_414)
            _1519 <= _5492;
        else
            _1519 <= _35;
    end
    assign _1556 = _1555 ? _1519 : _1539;
    assign _1552 = _1548 ? _1551 : _1539;
    assign _1557 = _1545 ? _1556 : _1552;
    assign _1558 = _1058 ? _1557 : _1539;
    assign _1544 = _1055 & _408;
    assign _1559 = _1544 ? _1551 : _1558;
    assign _36 = _1559;
    always @(posedge _416) begin
        if (_414)
            _1539 <= _5492;
        else
            _1539 <= _36;
    end
    assign _1565 = _1564 ? _1539 : _1551;
    assign _1573 = _1561 ? _1572 : _1565;
    assign _1574 = _1058 ? _1573 : _1551;
    assign _1560 = _1055 & _408;
    assign _1575 = _1560 ? _1571 : _1574;
    assign _37 = _1575;
    always @(posedge _416) begin
        if (_414)
            _1551 <= _5492;
        else
            _1551 <= _37;
    end
    assign _1588 = _1587 ? _1551 : _1571;
    assign _1584 = _1580 ? _1583 : _1571;
    assign _1589 = _1577 ? _1588 : _1584;
    assign _1590 = _1058 ? _1589 : _1571;
    assign _1576 = _1055 & _408;
    assign _1591 = _1576 ? _1583 : _1590;
    assign _38 = _1591;
    always @(posedge _416) begin
        if (_414)
            _1571 <= _5492;
        else
            _1571 <= _38;
    end
    assign _1597 = _1596 ? _1571 : _1583;
    assign _1605 = _1593 ? _1604 : _1597;
    assign _1606 = _1058 ? _1605 : _1583;
    assign _1592 = _1055 & _408;
    assign _1607 = _1592 ? _1603 : _1606;
    assign _39 = _1607;
    always @(posedge _416) begin
        if (_414)
            _1583 <= _5492;
        else
            _1583 <= _39;
    end
    assign _1620 = _1619 ? _1583 : _1603;
    assign _1616 = _1612 ? _1615 : _1603;
    assign _1621 = _1609 ? _1620 : _1616;
    assign _1622 = _1058 ? _1621 : _1603;
    assign _1608 = _1055 & _408;
    assign _1623 = _1608 ? _1615 : _1622;
    assign _40 = _1623;
    always @(posedge _416) begin
        if (_414)
            _1603 <= _5492;
        else
            _1603 <= _40;
    end
    assign _1629 = _1628 ? _1603 : _1615;
    assign _1637 = _1625 ? _1636 : _1629;
    assign _1638 = _1058 ? _1637 : _1615;
    assign _1624 = _1055 & _408;
    assign _1639 = _1624 ? _1635 : _1638;
    assign _41 = _1639;
    always @(posedge _416) begin
        if (_414)
            _1615 <= _5492;
        else
            _1615 <= _41;
    end
    assign _1652 = _1651 ? _1615 : _1635;
    assign _1648 = _1644 ? _1647 : _1635;
    assign _1653 = _1641 ? _1652 : _1648;
    assign _1654 = _1058 ? _1653 : _1635;
    assign _1640 = _1055 & _408;
    assign _1655 = _1640 ? _1647 : _1654;
    assign _42 = _1655;
    always @(posedge _416) begin
        if (_414)
            _1635 <= _5492;
        else
            _1635 <= _42;
    end
    assign _1661 = _1660 ? _1635 : _1647;
    assign _1669 = _1657 ? _1668 : _1661;
    assign _1670 = _1058 ? _1669 : _1647;
    assign _1656 = _1055 & _408;
    assign _1671 = _1656 ? _1667 : _1670;
    assign _43 = _1671;
    always @(posedge _416) begin
        if (_414)
            _1647 <= _5492;
        else
            _1647 <= _43;
    end
    assign _1684 = _1683 ? _1647 : _1667;
    assign _1680 = _1676 ? _1679 : _1667;
    assign _1685 = _1673 ? _1684 : _1680;
    assign _1686 = _1058 ? _1685 : _1667;
    assign _1672 = _1055 & _408;
    assign _1687 = _1672 ? _1679 : _1686;
    assign _44 = _1687;
    always @(posedge _416) begin
        if (_414)
            _1667 <= _5492;
        else
            _1667 <= _44;
    end
    assign _1693 = _1692 ? _1667 : _1679;
    assign _1701 = _1689 ? _1700 : _1693;
    assign _1702 = _1058 ? _1701 : _1679;
    assign _1688 = _1055 & _408;
    assign _1703 = _1688 ? _1699 : _1702;
    assign _45 = _1703;
    always @(posedge _416) begin
        if (_414)
            _1679 <= _5492;
        else
            _1679 <= _45;
    end
    assign _1716 = _1715 ? _1679 : _1699;
    assign _1712 = _1708 ? _1711 : _1699;
    assign _1717 = _1705 ? _1716 : _1712;
    assign _1718 = _1058 ? _1717 : _1699;
    assign _1704 = _1055 & _408;
    assign _1719 = _1704 ? _1711 : _1718;
    assign _46 = _1719;
    always @(posedge _416) begin
        if (_414)
            _1699 <= _5492;
        else
            _1699 <= _46;
    end
    assign _1725 = _1724 ? _1699 : _1711;
    assign _1733 = _1721 ? _1732 : _1725;
    assign _1734 = _1058 ? _1733 : _1711;
    assign _1720 = _1055 & _408;
    assign _1735 = _1720 ? _1731 : _1734;
    assign _47 = _1735;
    always @(posedge _416) begin
        if (_414)
            _1711 <= _5492;
        else
            _1711 <= _47;
    end
    assign _1748 = _1747 ? _1711 : _1731;
    assign _1744 = _1740 ? _1743 : _1731;
    assign _1749 = _1737 ? _1748 : _1744;
    assign _1750 = _1058 ? _1749 : _1731;
    assign _1736 = _1055 & _408;
    assign _1751 = _1736 ? _1743 : _1750;
    assign _48 = _1751;
    always @(posedge _416) begin
        if (_414)
            _1731 <= _5492;
        else
            _1731 <= _48;
    end
    assign _1757 = _1756 ? _1731 : _1743;
    assign _1765 = _1753 ? _1764 : _1757;
    assign _1766 = _1058 ? _1765 : _1743;
    assign _1752 = _1055 & _408;
    assign _1767 = _1752 ? _1763 : _1766;
    assign _49 = _1767;
    always @(posedge _416) begin
        if (_414)
            _1743 <= _5492;
        else
            _1743 <= _49;
    end
    assign _1780 = _1779 ? _1743 : _1763;
    assign _1776 = _1772 ? _1775 : _1763;
    assign _1781 = _1769 ? _1780 : _1776;
    assign _1782 = _1058 ? _1781 : _1763;
    assign _1768 = _1055 & _408;
    assign _1783 = _1768 ? _1775 : _1782;
    assign _50 = _1783;
    always @(posedge _416) begin
        if (_414)
            _1763 <= _5492;
        else
            _1763 <= _50;
    end
    assign _1789 = _1788 ? _1763 : _1775;
    assign _1797 = _1785 ? _1796 : _1789;
    assign _1798 = _1058 ? _1797 : _1775;
    assign _1784 = _1055 & _408;
    assign _1799 = _1784 ? _1795 : _1798;
    assign _51 = _1799;
    always @(posedge _416) begin
        if (_414)
            _1775 <= _5492;
        else
            _1775 <= _51;
    end
    assign _1812 = _1811 ? _1775 : _1795;
    assign _1808 = _1804 ? _1807 : _1795;
    assign _1813 = _1801 ? _1812 : _1808;
    assign _1814 = _1058 ? _1813 : _1795;
    assign _1800 = _1055 & _408;
    assign _1815 = _1800 ? _1807 : _1814;
    assign _52 = _1815;
    always @(posedge _416) begin
        if (_414)
            _1795 <= _5492;
        else
            _1795 <= _52;
    end
    assign _1821 = _1820 ? _1795 : _1807;
    assign _1829 = _1817 ? _1828 : _1821;
    assign _1830 = _1058 ? _1829 : _1807;
    assign _1816 = _1055 & _408;
    assign _1831 = _1816 ? _1827 : _1830;
    assign _53 = _1831;
    always @(posedge _416) begin
        if (_414)
            _1807 <= _5492;
        else
            _1807 <= _53;
    end
    assign _1844 = _1843 ? _1807 : _1827;
    assign _1840 = _1836 ? _1839 : _1827;
    assign _1845 = _1833 ? _1844 : _1840;
    assign _1846 = _1058 ? _1845 : _1827;
    assign _1832 = _1055 & _408;
    assign _1847 = _1832 ? _1839 : _1846;
    assign _54 = _1847;
    always @(posedge _416) begin
        if (_414)
            _1827 <= _5492;
        else
            _1827 <= _54;
    end
    assign _1853 = _1852 ? _1827 : _1839;
    assign _1861 = _1849 ? _1860 : _1853;
    assign _1862 = _1058 ? _1861 : _1839;
    assign _1848 = _1055 & _408;
    assign _1863 = _1848 ? _1859 : _1862;
    assign _55 = _1863;
    always @(posedge _416) begin
        if (_414)
            _1839 <= _5492;
        else
            _1839 <= _55;
    end
    assign _1876 = _1875 ? _1839 : _1859;
    assign _1872 = _1868 ? _1871 : _1859;
    assign _1877 = _1865 ? _1876 : _1872;
    assign _1878 = _1058 ? _1877 : _1859;
    assign _1864 = _1055 & _408;
    assign _1879 = _1864 ? _1871 : _1878;
    assign _56 = _1879;
    always @(posedge _416) begin
        if (_414)
            _1859 <= _5492;
        else
            _1859 <= _56;
    end
    assign _1885 = _1884 ? _1859 : _1871;
    assign _1893 = _1881 ? _1892 : _1885;
    assign _1894 = _1058 ? _1893 : _1871;
    assign _1880 = _1055 & _408;
    assign _1895 = _1880 ? _1891 : _1894;
    assign _57 = _1895;
    always @(posedge _416) begin
        if (_414)
            _1871 <= _5492;
        else
            _1871 <= _57;
    end
    assign _1908 = _1907 ? _1871 : _1891;
    assign _1904 = _1900 ? _1903 : _1891;
    assign _1909 = _1897 ? _1908 : _1904;
    assign _1910 = _1058 ? _1909 : _1891;
    assign _1896 = _1055 & _408;
    assign _1911 = _1896 ? _1903 : _1910;
    assign _58 = _1911;
    always @(posedge _416) begin
        if (_414)
            _1891 <= _5492;
        else
            _1891 <= _58;
    end
    assign _1917 = _1916 ? _1891 : _1903;
    assign _1925 = _1913 ? _1924 : _1917;
    assign _1926 = _1058 ? _1925 : _1903;
    assign _1912 = _1055 & _408;
    assign _1927 = _1912 ? _1923 : _1926;
    assign _59 = _1927;
    always @(posedge _416) begin
        if (_414)
            _1903 <= _5492;
        else
            _1903 <= _59;
    end
    assign _1940 = _1939 ? _1903 : _1923;
    assign _1936 = _1932 ? _1935 : _1923;
    assign _1941 = _1929 ? _1940 : _1936;
    assign _1942 = _1058 ? _1941 : _1923;
    assign _1928 = _1055 & _408;
    assign _1943 = _1928 ? _1935 : _1942;
    assign _60 = _1943;
    always @(posedge _416) begin
        if (_414)
            _1923 <= _5492;
        else
            _1923 <= _60;
    end
    assign _1949 = _1948 ? _1923 : _1935;
    assign _1957 = _1945 ? _1956 : _1949;
    assign _1958 = _1058 ? _1957 : _1935;
    assign _1944 = _1055 & _408;
    assign _1959 = _1944 ? _1955 : _1958;
    assign _61 = _1959;
    always @(posedge _416) begin
        if (_414)
            _1935 <= _5492;
        else
            _1935 <= _61;
    end
    assign _1972 = _1971 ? _1935 : _1955;
    assign _1968 = _1964 ? _1967 : _1955;
    assign _1973 = _1961 ? _1972 : _1968;
    assign _1974 = _1058 ? _1973 : _1955;
    assign _1960 = _1055 & _408;
    assign _1975 = _1960 ? _1967 : _1974;
    assign _62 = _1975;
    always @(posedge _416) begin
        if (_414)
            _1955 <= _5492;
        else
            _1955 <= _62;
    end
    assign _1981 = _1980 ? _1955 : _1967;
    assign _1989 = _1977 ? _1988 : _1981;
    assign _1990 = _1058 ? _1989 : _1967;
    assign _1976 = _1055 & _408;
    assign _1991 = _1976 ? _1987 : _1990;
    assign _63 = _1991;
    always @(posedge _416) begin
        if (_414)
            _1967 <= _5492;
        else
            _1967 <= _63;
    end
    assign _2004 = _2003 ? _1967 : _1987;
    assign _2000 = _1996 ? _1999 : _1987;
    assign _2005 = _1993 ? _2004 : _2000;
    assign _2006 = _1058 ? _2005 : _1987;
    assign _1992 = _1055 & _408;
    assign _2007 = _1992 ? _1999 : _2006;
    assign _64 = _2007;
    always @(posedge _416) begin
        if (_414)
            _1987 <= _5492;
        else
            _1987 <= _64;
    end
    assign _2013 = _2012 ? _1987 : _1999;
    assign _2021 = _2009 ? _2020 : _2013;
    assign _2022 = _1058 ? _2021 : _1999;
    assign _2008 = _1055 & _408;
    assign _2023 = _2008 ? _2019 : _2022;
    assign _65 = _2023;
    always @(posedge _416) begin
        if (_414)
            _1999 <= _5492;
        else
            _1999 <= _65;
    end
    assign _2036 = _2035 ? _1999 : _2019;
    assign _2032 = _2028 ? _2031 : _2019;
    assign _2037 = _2025 ? _2036 : _2032;
    assign _2038 = _1058 ? _2037 : _2019;
    assign _2024 = _1055 & _408;
    assign _2039 = _2024 ? _2031 : _2038;
    assign _66 = _2039;
    always @(posedge _416) begin
        if (_414)
            _2019 <= _5492;
        else
            _2019 <= _66;
    end
    assign _2045 = _2044 ? _2019 : _2031;
    assign _2053 = _2041 ? _2052 : _2045;
    assign _2054 = _1058 ? _2053 : _2031;
    assign _2040 = _1055 & _408;
    assign _2055 = _2040 ? _2051 : _2054;
    assign _67 = _2055;
    always @(posedge _416) begin
        if (_414)
            _2031 <= _5492;
        else
            _2031 <= _67;
    end
    assign _2068 = _2067 ? _2031 : _2051;
    assign _2064 = _2060 ? _2063 : _2051;
    assign _2069 = _2057 ? _2068 : _2064;
    assign _2070 = _1058 ? _2069 : _2051;
    assign _2056 = _1055 & _408;
    assign _2071 = _2056 ? _2063 : _2070;
    assign _68 = _2071;
    always @(posedge _416) begin
        if (_414)
            _2051 <= _5492;
        else
            _2051 <= _68;
    end
    assign _2077 = _2076 ? _2051 : _2063;
    assign _2085 = _2073 ? _2084 : _2077;
    assign _2086 = _1058 ? _2085 : _2063;
    assign _2072 = _1055 & _408;
    assign _2087 = _2072 ? _2083 : _2086;
    assign _69 = _2087;
    always @(posedge _416) begin
        if (_414)
            _2063 <= _5492;
        else
            _2063 <= _69;
    end
    assign _2100 = _2099 ? _2063 : _2083;
    assign _2096 = _2092 ? _2095 : _2083;
    assign _2101 = _2089 ? _2100 : _2096;
    assign _2102 = _1058 ? _2101 : _2083;
    assign _2088 = _1055 & _408;
    assign _2103 = _2088 ? _2095 : _2102;
    assign _70 = _2103;
    always @(posedge _416) begin
        if (_414)
            _2083 <= _5492;
        else
            _2083 <= _70;
    end
    assign _2109 = _2108 ? _2083 : _2095;
    assign _2117 = _2105 ? _2116 : _2109;
    assign _2118 = _1058 ? _2117 : _2095;
    assign _2104 = _1055 & _408;
    assign _2119 = _2104 ? _2115 : _2118;
    assign _71 = _2119;
    always @(posedge _416) begin
        if (_414)
            _2095 <= _5492;
        else
            _2095 <= _71;
    end
    assign _2132 = _2131 ? _2095 : _2115;
    assign _2128 = _2124 ? _2127 : _2115;
    assign _2133 = _2121 ? _2132 : _2128;
    assign _2134 = _1058 ? _2133 : _2115;
    assign _2120 = _1055 & _408;
    assign _2135 = _2120 ? _2127 : _2134;
    assign _72 = _2135;
    always @(posedge _416) begin
        if (_414)
            _2115 <= _5492;
        else
            _2115 <= _72;
    end
    assign _2141 = _2140 ? _2115 : _2127;
    assign _2149 = _2137 ? _2148 : _2141;
    assign _2150 = _1058 ? _2149 : _2127;
    assign _2136 = _1055 & _408;
    assign _2151 = _2136 ? _2147 : _2150;
    assign _73 = _2151;
    always @(posedge _416) begin
        if (_414)
            _2127 <= _5492;
        else
            _2127 <= _73;
    end
    assign _2164 = _2163 ? _2127 : _2147;
    assign _2160 = _2156 ? _2159 : _2147;
    assign _2165 = _2153 ? _2164 : _2160;
    assign _2166 = _1058 ? _2165 : _2147;
    assign _2152 = _1055 & _408;
    assign _2167 = _2152 ? _2159 : _2166;
    assign _74 = _2167;
    always @(posedge _416) begin
        if (_414)
            _2147 <= _5492;
        else
            _2147 <= _74;
    end
    assign _2173 = _2172 ? _2147 : _2159;
    assign _2181 = _2169 ? _2180 : _2173;
    assign _2182 = _1058 ? _2181 : _2159;
    assign _2168 = _1055 & _408;
    assign _2183 = _2168 ? _2179 : _2182;
    assign _75 = _2183;
    always @(posedge _416) begin
        if (_414)
            _2159 <= _5492;
        else
            _2159 <= _75;
    end
    assign _2196 = _2195 ? _2159 : _2179;
    assign _2192 = _2188 ? _2191 : _2179;
    assign _2197 = _2185 ? _2196 : _2192;
    assign _2198 = _1058 ? _2197 : _2179;
    assign _2184 = _1055 & _408;
    assign _2199 = _2184 ? _2191 : _2198;
    assign _76 = _2199;
    always @(posedge _416) begin
        if (_414)
            _2179 <= _5492;
        else
            _2179 <= _76;
    end
    assign _2205 = _2204 ? _2179 : _2191;
    assign _2213 = _2201 ? _2212 : _2205;
    assign _2214 = _1058 ? _2213 : _2191;
    assign _2200 = _1055 & _408;
    assign _2215 = _2200 ? _2211 : _2214;
    assign _77 = _2215;
    always @(posedge _416) begin
        if (_414)
            _2191 <= _5492;
        else
            _2191 <= _77;
    end
    assign _2228 = _2227 ? _2191 : _2211;
    assign _2224 = _2220 ? _2223 : _2211;
    assign _2229 = _2217 ? _2228 : _2224;
    assign _2230 = _1058 ? _2229 : _2211;
    assign _2216 = _1055 & _408;
    assign _2231 = _2216 ? _2223 : _2230;
    assign _78 = _2231;
    always @(posedge _416) begin
        if (_414)
            _2211 <= _5492;
        else
            _2211 <= _78;
    end
    assign _2237 = _2236 ? _2211 : _2223;
    assign _2245 = _2233 ? _2244 : _2237;
    assign _2246 = _1058 ? _2245 : _2223;
    assign _2232 = _1055 & _408;
    assign _2247 = _2232 ? _2243 : _2246;
    assign _79 = _2247;
    always @(posedge _416) begin
        if (_414)
            _2223 <= _5492;
        else
            _2223 <= _79;
    end
    assign _2260 = _2259 ? _2223 : _2243;
    assign _2256 = _2252 ? _2255 : _2243;
    assign _2261 = _2249 ? _2260 : _2256;
    assign _2262 = _1058 ? _2261 : _2243;
    assign _2248 = _1055 & _408;
    assign _2263 = _2248 ? _2255 : _2262;
    assign _80 = _2263;
    always @(posedge _416) begin
        if (_414)
            _2243 <= _5492;
        else
            _2243 <= _80;
    end
    assign _2269 = _2268 ? _2243 : _2255;
    assign _2277 = _2265 ? _2276 : _2269;
    assign _2278 = _1058 ? _2277 : _2255;
    assign _2264 = _1055 & _408;
    assign _2279 = _2264 ? _2275 : _2278;
    assign _81 = _2279;
    always @(posedge _416) begin
        if (_414)
            _2255 <= _5492;
        else
            _2255 <= _81;
    end
    assign _2292 = _2291 ? _2255 : _2275;
    assign _2288 = _2284 ? _2287 : _2275;
    assign _2293 = _2281 ? _2292 : _2288;
    assign _2294 = _1058 ? _2293 : _2275;
    assign _2280 = _1055 & _408;
    assign _2295 = _2280 ? _2287 : _2294;
    assign _82 = _2295;
    always @(posedge _416) begin
        if (_414)
            _2275 <= _5492;
        else
            _2275 <= _82;
    end
    assign _2301 = _2300 ? _2275 : _2287;
    assign _2309 = _2297 ? _2308 : _2301;
    assign _2310 = _1058 ? _2309 : _2287;
    assign _2296 = _1055 & _408;
    assign _2311 = _2296 ? _2307 : _2310;
    assign _83 = _2311;
    always @(posedge _416) begin
        if (_414)
            _2287 <= _5492;
        else
            _2287 <= _83;
    end
    assign _2324 = _2323 ? _2287 : _2307;
    assign _2320 = _2316 ? _2319 : _2307;
    assign _2325 = _2313 ? _2324 : _2320;
    assign _2326 = _1058 ? _2325 : _2307;
    assign _2312 = _1055 & _408;
    assign _2327 = _2312 ? _2319 : _2326;
    assign _84 = _2327;
    always @(posedge _416) begin
        if (_414)
            _2307 <= _5492;
        else
            _2307 <= _84;
    end
    assign _2333 = _2332 ? _2307 : _2319;
    assign _2341 = _2329 ? _2340 : _2333;
    assign _2342 = _1058 ? _2341 : _2319;
    assign _2328 = _1055 & _408;
    assign _2343 = _2328 ? _2339 : _2342;
    assign _85 = _2343;
    always @(posedge _416) begin
        if (_414)
            _2319 <= _5492;
        else
            _2319 <= _85;
    end
    assign _2356 = _2355 ? _2319 : _2339;
    assign _2352 = _2348 ? _2351 : _2339;
    assign _2357 = _2345 ? _2356 : _2352;
    assign _2358 = _1058 ? _2357 : _2339;
    assign _2344 = _1055 & _408;
    assign _2359 = _2344 ? _2351 : _2358;
    assign _86 = _2359;
    always @(posedge _416) begin
        if (_414)
            _2339 <= _5492;
        else
            _2339 <= _86;
    end
    assign _2365 = _2364 ? _2339 : _2351;
    assign _2373 = _2361 ? _2372 : _2365;
    assign _2374 = _1058 ? _2373 : _2351;
    assign _2360 = _1055 & _408;
    assign _2375 = _2360 ? _2371 : _2374;
    assign _87 = _2375;
    always @(posedge _416) begin
        if (_414)
            _2351 <= _5492;
        else
            _2351 <= _87;
    end
    assign _2388 = _2387 ? _2351 : _2371;
    assign _2384 = _2380 ? _2383 : _2371;
    assign _2389 = _2377 ? _2388 : _2384;
    assign _2390 = _1058 ? _2389 : _2371;
    assign _2376 = _1055 & _408;
    assign _2391 = _2376 ? _2383 : _2390;
    assign _88 = _2391;
    always @(posedge _416) begin
        if (_414)
            _2371 <= _5492;
        else
            _2371 <= _88;
    end
    assign _2397 = _2396 ? _2371 : _2383;
    assign _2405 = _2393 ? _2404 : _2397;
    assign _2406 = _1058 ? _2405 : _2383;
    assign _2392 = _1055 & _408;
    assign _2407 = _2392 ? _2403 : _2406;
    assign _89 = _2407;
    always @(posedge _416) begin
        if (_414)
            _2383 <= _5492;
        else
            _2383 <= _89;
    end
    assign _2420 = _2419 ? _2383 : _2403;
    assign _2416 = _2412 ? _2415 : _2403;
    assign _2421 = _2409 ? _2420 : _2416;
    assign _2422 = _1058 ? _2421 : _2403;
    assign _2408 = _1055 & _408;
    assign _2423 = _2408 ? _2415 : _2422;
    assign _90 = _2423;
    always @(posedge _416) begin
        if (_414)
            _2403 <= _5492;
        else
            _2403 <= _90;
    end
    assign _2429 = _2428 ? _2403 : _2415;
    assign _2437 = _2425 ? _2436 : _2429;
    assign _2438 = _1058 ? _2437 : _2415;
    assign _2424 = _1055 & _408;
    assign _2439 = _2424 ? _2435 : _2438;
    assign _91 = _2439;
    always @(posedge _416) begin
        if (_414)
            _2415 <= _5492;
        else
            _2415 <= _91;
    end
    assign _2452 = _2451 ? _2415 : _2435;
    assign _2448 = _2444 ? _2447 : _2435;
    assign _2453 = _2441 ? _2452 : _2448;
    assign _2454 = _1058 ? _2453 : _2435;
    assign _2440 = _1055 & _408;
    assign _2455 = _2440 ? _2447 : _2454;
    assign _92 = _2455;
    always @(posedge _416) begin
        if (_414)
            _2435 <= _5492;
        else
            _2435 <= _92;
    end
    assign _2461 = _2460 ? _2435 : _2447;
    assign _2469 = _2457 ? _2468 : _2461;
    assign _2470 = _1058 ? _2469 : _2447;
    assign _2456 = _1055 & _408;
    assign _2471 = _2456 ? _2467 : _2470;
    assign _93 = _2471;
    always @(posedge _416) begin
        if (_414)
            _2447 <= _5492;
        else
            _2447 <= _93;
    end
    assign _2484 = _2483 ? _2447 : _2467;
    assign _2480 = _2476 ? _2479 : _2467;
    assign _2485 = _2473 ? _2484 : _2480;
    assign _2486 = _1058 ? _2485 : _2467;
    assign _2472 = _1055 & _408;
    assign _2487 = _2472 ? _2479 : _2486;
    assign _94 = _2487;
    always @(posedge _416) begin
        if (_414)
            _2467 <= _5492;
        else
            _2467 <= _94;
    end
    assign _2493 = _2492 ? _2467 : _2479;
    assign _2501 = _2489 ? _2500 : _2493;
    assign _2502 = _1058 ? _2501 : _2479;
    assign _2488 = _1055 & _408;
    assign _2503 = _2488 ? _2499 : _2502;
    assign _95 = _2503;
    always @(posedge _416) begin
        if (_414)
            _2479 <= _5492;
        else
            _2479 <= _95;
    end
    assign _2516 = _2515 ? _2479 : _2499;
    assign _2512 = _2508 ? _2511 : _2499;
    assign _2517 = _2505 ? _2516 : _2512;
    assign _2518 = _1058 ? _2517 : _2499;
    assign _2504 = _1055 & _408;
    assign _2519 = _2504 ? _2511 : _2518;
    assign _96 = _2519;
    always @(posedge _416) begin
        if (_414)
            _2499 <= _5492;
        else
            _2499 <= _96;
    end
    assign _2525 = _2524 ? _2499 : _2511;
    assign _2533 = _2521 ? _2532 : _2525;
    assign _2534 = _1058 ? _2533 : _2511;
    assign _2520 = _1055 & _408;
    assign _2535 = _2520 ? _2531 : _2534;
    assign _97 = _2535;
    always @(posedge _416) begin
        if (_414)
            _2511 <= _5492;
        else
            _2511 <= _97;
    end
    assign _2548 = _2547 ? _2511 : _2531;
    assign _2544 = _2540 ? _2543 : _2531;
    assign _2549 = _2537 ? _2548 : _2544;
    assign _2550 = _1058 ? _2549 : _2531;
    assign _2536 = _1055 & _408;
    assign _2551 = _2536 ? _2543 : _2550;
    assign _98 = _2551;
    always @(posedge _416) begin
        if (_414)
            _2531 <= _5492;
        else
            _2531 <= _98;
    end
    assign _2557 = _2556 ? _2531 : _2543;
    assign _2565 = _2553 ? _2564 : _2557;
    assign _2566 = _1058 ? _2565 : _2543;
    assign _2552 = _1055 & _408;
    assign _2567 = _2552 ? _2563 : _2566;
    assign _99 = _2567;
    always @(posedge _416) begin
        if (_414)
            _2543 <= _5492;
        else
            _2543 <= _99;
    end
    assign _2580 = _2579 ? _2543 : _2563;
    assign _2576 = _2572 ? _2575 : _2563;
    assign _2581 = _2569 ? _2580 : _2576;
    assign _2582 = _1058 ? _2581 : _2563;
    assign _2568 = _1055 & _408;
    assign _2583 = _2568 ? _2575 : _2582;
    assign _100 = _2583;
    always @(posedge _416) begin
        if (_414)
            _2563 <= _5492;
        else
            _2563 <= _100;
    end
    assign _2589 = _2588 ? _2563 : _2575;
    assign _2597 = _2585 ? _2596 : _2589;
    assign _2598 = _1058 ? _2597 : _2575;
    assign _2584 = _1055 & _408;
    assign _2599 = _2584 ? _2595 : _2598;
    assign _101 = _2599;
    always @(posedge _416) begin
        if (_414)
            _2575 <= _5492;
        else
            _2575 <= _101;
    end
    assign _2612 = _2611 ? _2575 : _2595;
    assign _2608 = _2604 ? _2607 : _2595;
    assign _2613 = _2601 ? _2612 : _2608;
    assign _2614 = _1058 ? _2613 : _2595;
    assign _2600 = _1055 & _408;
    assign _2615 = _2600 ? _2607 : _2614;
    assign _102 = _2615;
    always @(posedge _416) begin
        if (_414)
            _2595 <= _5492;
        else
            _2595 <= _102;
    end
    assign _2621 = _2620 ? _2595 : _2607;
    assign _2629 = _2617 ? _2628 : _2621;
    assign _2630 = _1058 ? _2629 : _2607;
    assign _2616 = _1055 & _408;
    assign _2631 = _2616 ? _2627 : _2630;
    assign _103 = _2631;
    always @(posedge _416) begin
        if (_414)
            _2607 <= _5492;
        else
            _2607 <= _103;
    end
    assign _2644 = _2643 ? _2607 : _2627;
    assign _2640 = _2636 ? _2639 : _2627;
    assign _2645 = _2633 ? _2644 : _2640;
    assign _2646 = _1058 ? _2645 : _2627;
    assign _2632 = _1055 & _408;
    assign _2647 = _2632 ? _2639 : _2646;
    assign _104 = _2647;
    always @(posedge _416) begin
        if (_414)
            _2627 <= _5492;
        else
            _2627 <= _104;
    end
    assign _2653 = _2652 ? _2627 : _2639;
    assign _2661 = _2649 ? _2660 : _2653;
    assign _2662 = _1058 ? _2661 : _2639;
    assign _2648 = _1055 & _408;
    assign _2663 = _2648 ? _2659 : _2662;
    assign _105 = _2663;
    always @(posedge _416) begin
        if (_414)
            _2639 <= _5492;
        else
            _2639 <= _105;
    end
    assign _2676 = _2675 ? _2639 : _2659;
    assign _2672 = _2668 ? _2671 : _2659;
    assign _2677 = _2665 ? _2676 : _2672;
    assign _2678 = _1058 ? _2677 : _2659;
    assign _2664 = _1055 & _408;
    assign _2679 = _2664 ? _2671 : _2678;
    assign _106 = _2679;
    always @(posedge _416) begin
        if (_414)
            _2659 <= _5492;
        else
            _2659 <= _106;
    end
    assign _2685 = _2684 ? _2659 : _2671;
    assign _2693 = _2681 ? _2692 : _2685;
    assign _2694 = _1058 ? _2693 : _2671;
    assign _2680 = _1055 & _408;
    assign _2695 = _2680 ? _2691 : _2694;
    assign _107 = _2695;
    always @(posedge _416) begin
        if (_414)
            _2671 <= _5492;
        else
            _2671 <= _107;
    end
    assign _2708 = _2707 ? _2671 : _2691;
    assign _2704 = _2700 ? _2703 : _2691;
    assign _2709 = _2697 ? _2708 : _2704;
    assign _2710 = _1058 ? _2709 : _2691;
    assign _2696 = _1055 & _408;
    assign _2711 = _2696 ? _2703 : _2710;
    assign _108 = _2711;
    always @(posedge _416) begin
        if (_414)
            _2691 <= _5492;
        else
            _2691 <= _108;
    end
    assign _2717 = _2716 ? _2691 : _2703;
    assign _2725 = _2713 ? _2724 : _2717;
    assign _2726 = _1058 ? _2725 : _2703;
    assign _2712 = _1055 & _408;
    assign _2727 = _2712 ? _2723 : _2726;
    assign _109 = _2727;
    always @(posedge _416) begin
        if (_414)
            _2703 <= _5492;
        else
            _2703 <= _109;
    end
    assign _2740 = _2739 ? _2703 : _2723;
    assign _2736 = _2732 ? _2735 : _2723;
    assign _2741 = _2729 ? _2740 : _2736;
    assign _2742 = _1058 ? _2741 : _2723;
    assign _2728 = _1055 & _408;
    assign _2743 = _2728 ? _2735 : _2742;
    assign _110 = _2743;
    always @(posedge _416) begin
        if (_414)
            _2723 <= _5492;
        else
            _2723 <= _110;
    end
    assign _2749 = _2748 ? _2723 : _2735;
    assign _2757 = _2745 ? _2756 : _2749;
    assign _2758 = _1058 ? _2757 : _2735;
    assign _2744 = _1055 & _408;
    assign _2759 = _2744 ? _2755 : _2758;
    assign _111 = _2759;
    always @(posedge _416) begin
        if (_414)
            _2735 <= _5492;
        else
            _2735 <= _111;
    end
    assign _2772 = _2771 ? _2735 : _2755;
    assign _2768 = _2764 ? _2767 : _2755;
    assign _2773 = _2761 ? _2772 : _2768;
    assign _2774 = _1058 ? _2773 : _2755;
    assign _2760 = _1055 & _408;
    assign _2775 = _2760 ? _2767 : _2774;
    assign _112 = _2775;
    always @(posedge _416) begin
        if (_414)
            _2755 <= _5492;
        else
            _2755 <= _112;
    end
    assign _2781 = _2780 ? _2755 : _2767;
    assign _2789 = _2777 ? _2788 : _2781;
    assign _2790 = _1058 ? _2789 : _2767;
    assign _2776 = _1055 & _408;
    assign _2791 = _2776 ? _2787 : _2790;
    assign _113 = _2791;
    always @(posedge _416) begin
        if (_414)
            _2767 <= _5492;
        else
            _2767 <= _113;
    end
    assign _2804 = _2803 ? _2767 : _2787;
    assign _2800 = _2796 ? _2799 : _2787;
    assign _2805 = _2793 ? _2804 : _2800;
    assign _2806 = _1058 ? _2805 : _2787;
    assign _2792 = _1055 & _408;
    assign _2807 = _2792 ? _2799 : _2806;
    assign _114 = _2807;
    always @(posedge _416) begin
        if (_414)
            _2787 <= _5492;
        else
            _2787 <= _114;
    end
    assign _2813 = _2812 ? _2787 : _2799;
    assign _2821 = _2809 ? _2820 : _2813;
    assign _2822 = _1058 ? _2821 : _2799;
    assign _2808 = _1055 & _408;
    assign _2823 = _2808 ? _2819 : _2822;
    assign _115 = _2823;
    always @(posedge _416) begin
        if (_414)
            _2799 <= _5492;
        else
            _2799 <= _115;
    end
    assign _2836 = _2835 ? _2799 : _2819;
    assign _2832 = _2828 ? _2831 : _2819;
    assign _2837 = _2825 ? _2836 : _2832;
    assign _2838 = _1058 ? _2837 : _2819;
    assign _2824 = _1055 & _408;
    assign _2839 = _2824 ? _2831 : _2838;
    assign _116 = _2839;
    always @(posedge _416) begin
        if (_414)
            _2819 <= _5492;
        else
            _2819 <= _116;
    end
    assign _2845 = _2844 ? _2819 : _2831;
    assign _2853 = _2841 ? _2852 : _2845;
    assign _2854 = _1058 ? _2853 : _2831;
    assign _2840 = _1055 & _408;
    assign _2855 = _2840 ? _2851 : _2854;
    assign _117 = _2855;
    always @(posedge _416) begin
        if (_414)
            _2831 <= _5492;
        else
            _2831 <= _117;
    end
    assign _2868 = _2867 ? _2831 : _2851;
    assign _2864 = _2860 ? _2863 : _2851;
    assign _2869 = _2857 ? _2868 : _2864;
    assign _2870 = _1058 ? _2869 : _2851;
    assign _2856 = _1055 & _408;
    assign _2871 = _2856 ? _2863 : _2870;
    assign _118 = _2871;
    always @(posedge _416) begin
        if (_414)
            _2851 <= _5492;
        else
            _2851 <= _118;
    end
    assign _2877 = _2876 ? _2851 : _2863;
    assign _2885 = _2873 ? _2884 : _2877;
    assign _2886 = _1058 ? _2885 : _2863;
    assign _2872 = _1055 & _408;
    assign _2887 = _2872 ? _2883 : _2886;
    assign _119 = _2887;
    always @(posedge _416) begin
        if (_414)
            _2863 <= _5492;
        else
            _2863 <= _119;
    end
    assign _2900 = _2899 ? _2863 : _2883;
    assign _2896 = _2892 ? _2895 : _2883;
    assign _2901 = _2889 ? _2900 : _2896;
    assign _2902 = _1058 ? _2901 : _2883;
    assign _2888 = _1055 & _408;
    assign _2903 = _2888 ? _2895 : _2902;
    assign _120 = _2903;
    always @(posedge _416) begin
        if (_414)
            _2883 <= _5492;
        else
            _2883 <= _120;
    end
    assign _2909 = _2908 ? _2883 : _2895;
    assign _2917 = _2905 ? _2916 : _2909;
    assign _2918 = _1058 ? _2917 : _2895;
    assign _2904 = _1055 & _408;
    assign _2919 = _2904 ? _2915 : _2918;
    assign _121 = _2919;
    always @(posedge _416) begin
        if (_414)
            _2895 <= _5492;
        else
            _2895 <= _121;
    end
    assign _2932 = _2931 ? _2895 : _2915;
    assign _2928 = _2924 ? _2927 : _2915;
    assign _2933 = _2921 ? _2932 : _2928;
    assign _2934 = _1058 ? _2933 : _2915;
    assign _2920 = _1055 & _408;
    assign _2935 = _2920 ? _2927 : _2934;
    assign _122 = _2935;
    always @(posedge _416) begin
        if (_414)
            _2915 <= _5492;
        else
            _2915 <= _122;
    end
    assign _2941 = _2940 ? _2915 : _2927;
    assign _2949 = _2937 ? _2948 : _2941;
    assign _2950 = _1058 ? _2949 : _2927;
    assign _2936 = _1055 & _408;
    assign _2951 = _2936 ? _2947 : _2950;
    assign _123 = _2951;
    always @(posedge _416) begin
        if (_414)
            _2927 <= _5492;
        else
            _2927 <= _123;
    end
    assign _2964 = _2963 ? _2927 : _2947;
    assign _2960 = _2956 ? _2959 : _2947;
    assign _2965 = _2953 ? _2964 : _2960;
    assign _2966 = _1058 ? _2965 : _2947;
    assign _2952 = _1055 & _408;
    assign _2967 = _2952 ? _2959 : _2966;
    assign _124 = _2967;
    always @(posedge _416) begin
        if (_414)
            _2947 <= _5492;
        else
            _2947 <= _124;
    end
    assign _2973 = _2972 ? _2947 : _2959;
    assign _2981 = _2969 ? _2980 : _2973;
    assign _2982 = _1058 ? _2981 : _2959;
    assign _2968 = _1055 & _408;
    assign _2983 = _2968 ? _2979 : _2982;
    assign _125 = _2983;
    always @(posedge _416) begin
        if (_414)
            _2959 <= _5492;
        else
            _2959 <= _125;
    end
    assign _2996 = _2995 ? _2959 : _2979;
    assign _2992 = _2988 ? _2991 : _2979;
    assign _2997 = _2985 ? _2996 : _2992;
    assign _2998 = _1058 ? _2997 : _2979;
    assign _2984 = _1055 & _408;
    assign _2999 = _2984 ? _2991 : _2998;
    assign _126 = _2999;
    always @(posedge _416) begin
        if (_414)
            _2979 <= _5492;
        else
            _2979 <= _126;
    end
    assign _3005 = _3004 ? _2979 : _2991;
    assign _3013 = _3001 ? _3012 : _3005;
    assign _3014 = _1058 ? _3013 : _2991;
    assign _3000 = _1055 & _408;
    assign _3015 = _3000 ? _3011 : _3014;
    assign _127 = _3015;
    always @(posedge _416) begin
        if (_414)
            _2991 <= _5492;
        else
            _2991 <= _127;
    end
    assign _3028 = _3027 ? _2991 : _3011;
    assign _3024 = _3020 ? _3023 : _3011;
    assign _3029 = _3017 ? _3028 : _3024;
    assign _3030 = _1058 ? _3029 : _3011;
    assign _3016 = _1055 & _408;
    assign _3031 = _3016 ? _3023 : _3030;
    assign _128 = _3031;
    always @(posedge _416) begin
        if (_414)
            _3011 <= _5492;
        else
            _3011 <= _128;
    end
    assign _3037 = _3036 ? _3011 : _3023;
    assign _3045 = _3033 ? _3044 : _3037;
    assign _3046 = _1058 ? _3045 : _3023;
    assign _3032 = _1055 & _408;
    assign _3047 = _3032 ? _3043 : _3046;
    assign _129 = _3047;
    always @(posedge _416) begin
        if (_414)
            _3023 <= _5492;
        else
            _3023 <= _129;
    end
    assign _3060 = _3059 ? _3023 : _3043;
    assign _3056 = _3052 ? _3055 : _3043;
    assign _3061 = _3049 ? _3060 : _3056;
    assign _3062 = _1058 ? _3061 : _3043;
    assign _3048 = _1055 & _408;
    assign _3063 = _3048 ? _3055 : _3062;
    assign _130 = _3063;
    always @(posedge _416) begin
        if (_414)
            _3043 <= _5492;
        else
            _3043 <= _130;
    end
    assign _3069 = _3068 ? _3043 : _3055;
    assign _3077 = _3065 ? _3076 : _3069;
    assign _3078 = _1058 ? _3077 : _3055;
    assign _3064 = _1055 & _408;
    assign _3079 = _3064 ? _3075 : _3078;
    assign _131 = _3079;
    always @(posedge _416) begin
        if (_414)
            _3055 <= _5492;
        else
            _3055 <= _131;
    end
    assign _3092 = _3091 ? _3055 : _3075;
    assign _3088 = _3084 ? _3087 : _3075;
    assign _3093 = _3081 ? _3092 : _3088;
    assign _3094 = _1058 ? _3093 : _3075;
    assign _3080 = _1055 & _408;
    assign _3095 = _3080 ? _3087 : _3094;
    assign _132 = _3095;
    always @(posedge _416) begin
        if (_414)
            _3075 <= _5492;
        else
            _3075 <= _132;
    end
    assign _3101 = _3100 ? _3075 : _3087;
    assign _3109 = _3097 ? _3108 : _3101;
    assign _3110 = _1058 ? _3109 : _3087;
    assign _3096 = _1055 & _408;
    assign _3111 = _3096 ? _3107 : _3110;
    assign _133 = _3111;
    always @(posedge _416) begin
        if (_414)
            _3087 <= _5492;
        else
            _3087 <= _133;
    end
    assign _3124 = _3123 ? _3087 : _3107;
    assign _3120 = _3116 ? _3119 : _3107;
    assign _3125 = _3113 ? _3124 : _3120;
    assign _3126 = _1058 ? _3125 : _3107;
    assign _3112 = _1055 & _408;
    assign _3127 = _3112 ? _3119 : _3126;
    assign _134 = _3127;
    always @(posedge _416) begin
        if (_414)
            _3107 <= _5492;
        else
            _3107 <= _134;
    end
    assign _3133 = _3132 ? _3107 : _3119;
    assign _3141 = _3129 ? _3140 : _3133;
    assign _3142 = _1058 ? _3141 : _3119;
    assign _3128 = _1055 & _408;
    assign _3143 = _3128 ? _3139 : _3142;
    assign _135 = _3143;
    always @(posedge _416) begin
        if (_414)
            _3119 <= _5492;
        else
            _3119 <= _135;
    end
    assign _3156 = _3155 ? _3119 : _3139;
    assign _3152 = _3148 ? _3151 : _3139;
    assign _3157 = _3145 ? _3156 : _3152;
    assign _3158 = _1058 ? _3157 : _3139;
    assign _3144 = _1055 & _408;
    assign _3159 = _3144 ? _3151 : _3158;
    assign _136 = _3159;
    always @(posedge _416) begin
        if (_414)
            _3139 <= _5492;
        else
            _3139 <= _136;
    end
    assign _3165 = _3164 ? _3139 : _3151;
    assign _3173 = _3161 ? _3172 : _3165;
    assign _3174 = _1058 ? _3173 : _3151;
    assign _3160 = _1055 & _408;
    assign _3175 = _3160 ? _3171 : _3174;
    assign _137 = _3175;
    always @(posedge _416) begin
        if (_414)
            _3151 <= _5492;
        else
            _3151 <= _137;
    end
    assign _3188 = _3187 ? _3151 : _3171;
    assign _3184 = _3180 ? _3183 : _3171;
    assign _3189 = _3177 ? _3188 : _3184;
    assign _3190 = _1058 ? _3189 : _3171;
    assign _3176 = _1055 & _408;
    assign _3191 = _3176 ? _3183 : _3190;
    assign _138 = _3191;
    always @(posedge _416) begin
        if (_414)
            _3171 <= _5492;
        else
            _3171 <= _138;
    end
    assign _3197 = _3196 ? _3171 : _3183;
    assign _3205 = _3193 ? _3204 : _3197;
    assign _3206 = _1058 ? _3205 : _3183;
    assign _3192 = _1055 & _408;
    assign _3207 = _3192 ? _3203 : _3206;
    assign _139 = _3207;
    always @(posedge _416) begin
        if (_414)
            _3183 <= _5492;
        else
            _3183 <= _139;
    end
    assign _3220 = _3219 ? _3183 : _3203;
    assign _3216 = _3212 ? _3215 : _3203;
    assign _3221 = _3209 ? _3220 : _3216;
    assign _3222 = _1058 ? _3221 : _3203;
    assign _3208 = _1055 & _408;
    assign _3223 = _3208 ? _3215 : _3222;
    assign _140 = _3223;
    always @(posedge _416) begin
        if (_414)
            _3203 <= _5492;
        else
            _3203 <= _140;
    end
    assign _3229 = _3228 ? _3203 : _3215;
    assign _3237 = _3225 ? _3236 : _3229;
    assign _3238 = _1058 ? _3237 : _3215;
    assign _3224 = _1055 & _408;
    assign _3239 = _3224 ? _3235 : _3238;
    assign _141 = _3239;
    always @(posedge _416) begin
        if (_414)
            _3215 <= _5492;
        else
            _3215 <= _141;
    end
    assign _3252 = _3251 ? _3215 : _3235;
    assign _3248 = _3244 ? _3247 : _3235;
    assign _3253 = _3241 ? _3252 : _3248;
    assign _3254 = _1058 ? _3253 : _3235;
    assign _3240 = _1055 & _408;
    assign _3255 = _3240 ? _3247 : _3254;
    assign _142 = _3255;
    always @(posedge _416) begin
        if (_414)
            _3235 <= _5492;
        else
            _3235 <= _142;
    end
    assign _3261 = _3260 ? _3235 : _3247;
    assign _3269 = _3257 ? _3268 : _3261;
    assign _3270 = _1058 ? _3269 : _3247;
    assign _3256 = _1055 & _408;
    assign _3271 = _3256 ? _3267 : _3270;
    assign _143 = _3271;
    always @(posedge _416) begin
        if (_414)
            _3247 <= _5492;
        else
            _3247 <= _143;
    end
    assign _3284 = _3283 ? _3247 : _3267;
    assign _3280 = _3276 ? _3279 : _3267;
    assign _3285 = _3273 ? _3284 : _3280;
    assign _3286 = _1058 ? _3285 : _3267;
    assign _3272 = _1055 & _408;
    assign _3287 = _3272 ? _3279 : _3286;
    assign _144 = _3287;
    always @(posedge _416) begin
        if (_414)
            _3267 <= _5492;
        else
            _3267 <= _144;
    end
    assign _3293 = _3292 ? _3267 : _3279;
    assign _3301 = _3289 ? _3300 : _3293;
    assign _3302 = _1058 ? _3301 : _3279;
    assign _3288 = _1055 & _408;
    assign _3303 = _3288 ? _3299 : _3302;
    assign _145 = _3303;
    always @(posedge _416) begin
        if (_414)
            _3279 <= _5492;
        else
            _3279 <= _145;
    end
    assign _3316 = _3315 ? _3279 : _3299;
    assign _3312 = _3308 ? _3311 : _3299;
    assign _3317 = _3305 ? _3316 : _3312;
    assign _3318 = _1058 ? _3317 : _3299;
    assign _3304 = _1055 & _408;
    assign _3319 = _3304 ? _3311 : _3318;
    assign _146 = _3319;
    always @(posedge _416) begin
        if (_414)
            _3299 <= _5492;
        else
            _3299 <= _146;
    end
    assign _3325 = _3324 ? _3299 : _3311;
    assign _3333 = _3321 ? _3332 : _3325;
    assign _3334 = _1058 ? _3333 : _3311;
    assign _3320 = _1055 & _408;
    assign _3335 = _3320 ? _3331 : _3334;
    assign _147 = _3335;
    always @(posedge _416) begin
        if (_414)
            _3311 <= _5492;
        else
            _3311 <= _147;
    end
    assign _3348 = _3347 ? _3311 : _3331;
    assign _3344 = _3340 ? _3343 : _3331;
    assign _3349 = _3337 ? _3348 : _3344;
    assign _3350 = _1058 ? _3349 : _3331;
    assign _3336 = _1055 & _408;
    assign _3351 = _3336 ? _3343 : _3350;
    assign _148 = _3351;
    always @(posedge _416) begin
        if (_414)
            _3331 <= _5492;
        else
            _3331 <= _148;
    end
    assign _3357 = _3356 ? _3331 : _3343;
    assign _3365 = _3353 ? _3364 : _3357;
    assign _3366 = _1058 ? _3365 : _3343;
    assign _3352 = _1055 & _408;
    assign _3367 = _3352 ? _3363 : _3366;
    assign _149 = _3367;
    always @(posedge _416) begin
        if (_414)
            _3343 <= _5492;
        else
            _3343 <= _149;
    end
    assign _3380 = _3379 ? _3343 : _3363;
    assign _3376 = _3372 ? _3375 : _3363;
    assign _3381 = _3369 ? _3380 : _3376;
    assign _3382 = _1058 ? _3381 : _3363;
    assign _3368 = _1055 & _408;
    assign _3383 = _3368 ? _3375 : _3382;
    assign _150 = _3383;
    always @(posedge _416) begin
        if (_414)
            _3363 <= _5492;
        else
            _3363 <= _150;
    end
    assign _3389 = _3388 ? _3363 : _3375;
    assign _3397 = _3385 ? _3396 : _3389;
    assign _3398 = _1058 ? _3397 : _3375;
    assign _3384 = _1055 & _408;
    assign _3399 = _3384 ? _3395 : _3398;
    assign _151 = _3399;
    always @(posedge _416) begin
        if (_414)
            _3375 <= _5492;
        else
            _3375 <= _151;
    end
    assign _3412 = _3411 ? _3375 : _3395;
    assign _3408 = _3404 ? _3407 : _3395;
    assign _3413 = _3401 ? _3412 : _3408;
    assign _3414 = _1058 ? _3413 : _3395;
    assign _3400 = _1055 & _408;
    assign _3415 = _3400 ? _3407 : _3414;
    assign _152 = _3415;
    always @(posedge _416) begin
        if (_414)
            _3395 <= _5492;
        else
            _3395 <= _152;
    end
    assign _3421 = _3420 ? _3395 : _3407;
    assign _3429 = _3417 ? _3428 : _3421;
    assign _3430 = _1058 ? _3429 : _3407;
    assign _3416 = _1055 & _408;
    assign _3431 = _3416 ? _3427 : _3430;
    assign _153 = _3431;
    always @(posedge _416) begin
        if (_414)
            _3407 <= _5492;
        else
            _3407 <= _153;
    end
    assign _3444 = _3443 ? _3407 : _3427;
    assign _3440 = _3436 ? _3439 : _3427;
    assign _3445 = _3433 ? _3444 : _3440;
    assign _3446 = _1058 ? _3445 : _3427;
    assign _3432 = _1055 & _408;
    assign _3447 = _3432 ? _3439 : _3446;
    assign _154 = _3447;
    always @(posedge _416) begin
        if (_414)
            _3427 <= _5492;
        else
            _3427 <= _154;
    end
    assign _3453 = _3452 ? _3427 : _3439;
    assign _3461 = _3449 ? _3460 : _3453;
    assign _3462 = _1058 ? _3461 : _3439;
    assign _3448 = _1055 & _408;
    assign _3463 = _3448 ? _3459 : _3462;
    assign _155 = _3463;
    always @(posedge _416) begin
        if (_414)
            _3439 <= _5492;
        else
            _3439 <= _155;
    end
    assign _3476 = _3475 ? _3439 : _3459;
    assign _3472 = _3468 ? _3471 : _3459;
    assign _3477 = _3465 ? _3476 : _3472;
    assign _3478 = _1058 ? _3477 : _3459;
    assign _3464 = _1055 & _408;
    assign _3479 = _3464 ? _3471 : _3478;
    assign _156 = _3479;
    always @(posedge _416) begin
        if (_414)
            _3459 <= _5492;
        else
            _3459 <= _156;
    end
    assign _3485 = _3484 ? _3459 : _3471;
    assign _3493 = _3481 ? _3492 : _3485;
    assign _3494 = _1058 ? _3493 : _3471;
    assign _3480 = _1055 & _408;
    assign _3495 = _3480 ? _3491 : _3494;
    assign _157 = _3495;
    always @(posedge _416) begin
        if (_414)
            _3471 <= _5492;
        else
            _3471 <= _157;
    end
    assign _3508 = _3507 ? _3471 : _3491;
    assign _3504 = _3500 ? _3503 : _3491;
    assign _3509 = _3497 ? _3508 : _3504;
    assign _3510 = _1058 ? _3509 : _3491;
    assign _3496 = _1055 & _408;
    assign _3511 = _3496 ? _3503 : _3510;
    assign _158 = _3511;
    always @(posedge _416) begin
        if (_414)
            _3491 <= _5492;
        else
            _3491 <= _158;
    end
    assign _3517 = _3516 ? _3491 : _3503;
    assign _3525 = _3513 ? _3524 : _3517;
    assign _3526 = _1058 ? _3525 : _3503;
    assign _3512 = _1055 & _408;
    assign _3527 = _3512 ? _3523 : _3526;
    assign _159 = _3527;
    always @(posedge _416) begin
        if (_414)
            _3503 <= _5492;
        else
            _3503 <= _159;
    end
    assign _3540 = _3539 ? _3503 : _3523;
    assign _3536 = _3532 ? _3535 : _3523;
    assign _3541 = _3529 ? _3540 : _3536;
    assign _3542 = _1058 ? _3541 : _3523;
    assign _3528 = _1055 & _408;
    assign _3543 = _3528 ? _3535 : _3542;
    assign _160 = _3543;
    always @(posedge _416) begin
        if (_414)
            _3523 <= _5492;
        else
            _3523 <= _160;
    end
    assign _3549 = _3548 ? _3523 : _3535;
    assign _3557 = _3545 ? _3556 : _3549;
    assign _3558 = _1058 ? _3557 : _3535;
    assign _3544 = _1055 & _408;
    assign _3559 = _3544 ? _3555 : _3558;
    assign _161 = _3559;
    always @(posedge _416) begin
        if (_414)
            _3535 <= _5492;
        else
            _3535 <= _161;
    end
    assign _3572 = _3571 ? _3535 : _3555;
    assign _3568 = _3564 ? _3567 : _3555;
    assign _3573 = _3561 ? _3572 : _3568;
    assign _3574 = _1058 ? _3573 : _3555;
    assign _3560 = _1055 & _408;
    assign _3575 = _3560 ? _3567 : _3574;
    assign _162 = _3575;
    always @(posedge _416) begin
        if (_414)
            _3555 <= _5492;
        else
            _3555 <= _162;
    end
    assign _3581 = _3580 ? _3555 : _3567;
    assign _3589 = _3577 ? _3588 : _3581;
    assign _3590 = _1058 ? _3589 : _3567;
    assign _3576 = _1055 & _408;
    assign _3591 = _3576 ? _3587 : _3590;
    assign _163 = _3591;
    always @(posedge _416) begin
        if (_414)
            _3567 <= _5492;
        else
            _3567 <= _163;
    end
    assign _3604 = _3603 ? _3567 : _3587;
    assign _3600 = _3596 ? _3599 : _3587;
    assign _3605 = _3593 ? _3604 : _3600;
    assign _3606 = _1058 ? _3605 : _3587;
    assign _3592 = _1055 & _408;
    assign _3607 = _3592 ? _3599 : _3606;
    assign _164 = _3607;
    always @(posedge _416) begin
        if (_414)
            _3587 <= _5492;
        else
            _3587 <= _164;
    end
    assign _3613 = _3612 ? _3587 : _3599;
    assign _3621 = _3609 ? _3620 : _3613;
    assign _3622 = _1058 ? _3621 : _3599;
    assign _3608 = _1055 & _408;
    assign _3623 = _3608 ? _3619 : _3622;
    assign _165 = _3623;
    always @(posedge _416) begin
        if (_414)
            _3599 <= _5492;
        else
            _3599 <= _165;
    end
    assign _3636 = _3635 ? _3599 : _3619;
    assign _3632 = _3628 ? _3631 : _3619;
    assign _3637 = _3625 ? _3636 : _3632;
    assign _3638 = _1058 ? _3637 : _3619;
    assign _3624 = _1055 & _408;
    assign _3639 = _3624 ? _3631 : _3638;
    assign _166 = _3639;
    always @(posedge _416) begin
        if (_414)
            _3619 <= _5492;
        else
            _3619 <= _166;
    end
    assign _3645 = _3644 ? _3619 : _3631;
    assign _3653 = _3641 ? _3652 : _3645;
    assign _3654 = _1058 ? _3653 : _3631;
    assign _3640 = _1055 & _408;
    assign _3655 = _3640 ? _3651 : _3654;
    assign _167 = _3655;
    always @(posedge _416) begin
        if (_414)
            _3631 <= _5492;
        else
            _3631 <= _167;
    end
    assign _3668 = _3667 ? _3631 : _3651;
    assign _3664 = _3660 ? _3663 : _3651;
    assign _3669 = _3657 ? _3668 : _3664;
    assign _3670 = _1058 ? _3669 : _3651;
    assign _3656 = _1055 & _408;
    assign _3671 = _3656 ? _3663 : _3670;
    assign _168 = _3671;
    always @(posedge _416) begin
        if (_414)
            _3651 <= _5492;
        else
            _3651 <= _168;
    end
    assign _3677 = _3676 ? _3651 : _3663;
    assign _3685 = _3673 ? _3684 : _3677;
    assign _3686 = _1058 ? _3685 : _3663;
    assign _3672 = _1055 & _408;
    assign _3687 = _3672 ? _3683 : _3686;
    assign _169 = _3687;
    always @(posedge _416) begin
        if (_414)
            _3663 <= _5492;
        else
            _3663 <= _169;
    end
    assign _3700 = _3699 ? _3663 : _3683;
    assign _3696 = _3692 ? _3695 : _3683;
    assign _3701 = _3689 ? _3700 : _3696;
    assign _3702 = _1058 ? _3701 : _3683;
    assign _3688 = _1055 & _408;
    assign _3703 = _3688 ? _3695 : _3702;
    assign _170 = _3703;
    always @(posedge _416) begin
        if (_414)
            _3683 <= _5492;
        else
            _3683 <= _170;
    end
    assign _3709 = _3708 ? _3683 : _3695;
    assign _3717 = _3705 ? _3716 : _3709;
    assign _3718 = _1058 ? _3717 : _3695;
    assign _3704 = _1055 & _408;
    assign _3719 = _3704 ? _3715 : _3718;
    assign _171 = _3719;
    always @(posedge _416) begin
        if (_414)
            _3695 <= _5492;
        else
            _3695 <= _171;
    end
    assign _3732 = _3731 ? _3695 : _3715;
    assign _3728 = _3724 ? _3727 : _3715;
    assign _3733 = _3721 ? _3732 : _3728;
    assign _3734 = _1058 ? _3733 : _3715;
    assign _3720 = _1055 & _408;
    assign _3735 = _3720 ? _3727 : _3734;
    assign _172 = _3735;
    always @(posedge _416) begin
        if (_414)
            _3715 <= _5492;
        else
            _3715 <= _172;
    end
    assign _3741 = _3740 ? _3715 : _3727;
    assign _3749 = _3737 ? _3748 : _3741;
    assign _3750 = _1058 ? _3749 : _3727;
    assign _3736 = _1055 & _408;
    assign _3751 = _3736 ? _3747 : _3750;
    assign _173 = _3751;
    always @(posedge _416) begin
        if (_414)
            _3727 <= _5492;
        else
            _3727 <= _173;
    end
    assign _3764 = _3763 ? _3727 : _3747;
    assign _3760 = _3756 ? _3759 : _3747;
    assign _3765 = _3753 ? _3764 : _3760;
    assign _3766 = _1058 ? _3765 : _3747;
    assign _3752 = _1055 & _408;
    assign _3767 = _3752 ? _3759 : _3766;
    assign _174 = _3767;
    always @(posedge _416) begin
        if (_414)
            _3747 <= _5492;
        else
            _3747 <= _174;
    end
    assign _3773 = _3772 ? _3747 : _3759;
    assign _3781 = _3769 ? _3780 : _3773;
    assign _3782 = _1058 ? _3781 : _3759;
    assign _3768 = _1055 & _408;
    assign _3783 = _3768 ? _3779 : _3782;
    assign _175 = _3783;
    always @(posedge _416) begin
        if (_414)
            _3759 <= _5492;
        else
            _3759 <= _175;
    end
    assign _3796 = _3795 ? _3759 : _3779;
    assign _3792 = _3788 ? _3791 : _3779;
    assign _3797 = _3785 ? _3796 : _3792;
    assign _3798 = _1058 ? _3797 : _3779;
    assign _3784 = _1055 & _408;
    assign _3799 = _3784 ? _3791 : _3798;
    assign _176 = _3799;
    always @(posedge _416) begin
        if (_414)
            _3779 <= _5492;
        else
            _3779 <= _176;
    end
    assign _3805 = _3804 ? _3779 : _3791;
    assign _3813 = _3801 ? _3812 : _3805;
    assign _3814 = _1058 ? _3813 : _3791;
    assign _3800 = _1055 & _408;
    assign _3815 = _3800 ? _3811 : _3814;
    assign _177 = _3815;
    always @(posedge _416) begin
        if (_414)
            _3791 <= _5492;
        else
            _3791 <= _177;
    end
    assign _3828 = _3827 ? _3791 : _3811;
    assign _3824 = _3820 ? _3823 : _3811;
    assign _3829 = _3817 ? _3828 : _3824;
    assign _3830 = _1058 ? _3829 : _3811;
    assign _3816 = _1055 & _408;
    assign _3831 = _3816 ? _3823 : _3830;
    assign _178 = _3831;
    always @(posedge _416) begin
        if (_414)
            _3811 <= _5492;
        else
            _3811 <= _178;
    end
    assign _3837 = _3836 ? _3811 : _3823;
    assign _3845 = _3833 ? _3844 : _3837;
    assign _3846 = _1058 ? _3845 : _3823;
    assign _3832 = _1055 & _408;
    assign _3847 = _3832 ? _3843 : _3846;
    assign _179 = _3847;
    always @(posedge _416) begin
        if (_414)
            _3823 <= _5492;
        else
            _3823 <= _179;
    end
    assign _3860 = _3859 ? _3823 : _3843;
    assign _3856 = _3852 ? _3855 : _3843;
    assign _3861 = _3849 ? _3860 : _3856;
    assign _3862 = _1058 ? _3861 : _3843;
    assign _3848 = _1055 & _408;
    assign _3863 = _3848 ? _3855 : _3862;
    assign _180 = _3863;
    always @(posedge _416) begin
        if (_414)
            _3843 <= _5492;
        else
            _3843 <= _180;
    end
    assign _3869 = _3868 ? _3843 : _3855;
    assign _3877 = _3865 ? _3876 : _3869;
    assign _3878 = _1058 ? _3877 : _3855;
    assign _3864 = _1055 & _408;
    assign _3879 = _3864 ? _3875 : _3878;
    assign _181 = _3879;
    always @(posedge _416) begin
        if (_414)
            _3855 <= _5492;
        else
            _3855 <= _181;
    end
    assign _3892 = _3891 ? _3855 : _3875;
    assign _3888 = _3884 ? _3887 : _3875;
    assign _3893 = _3881 ? _3892 : _3888;
    assign _3894 = _1058 ? _3893 : _3875;
    assign _3880 = _1055 & _408;
    assign _3895 = _3880 ? _3887 : _3894;
    assign _182 = _3895;
    always @(posedge _416) begin
        if (_414)
            _3875 <= _5492;
        else
            _3875 <= _182;
    end
    assign _3901 = _3900 ? _3875 : _3887;
    assign _3909 = _3897 ? _3908 : _3901;
    assign _3910 = _1058 ? _3909 : _3887;
    assign _3896 = _1055 & _408;
    assign _3911 = _3896 ? _3907 : _3910;
    assign _183 = _3911;
    always @(posedge _416) begin
        if (_414)
            _3887 <= _5492;
        else
            _3887 <= _183;
    end
    assign _3924 = _3923 ? _3887 : _3907;
    assign _3920 = _3916 ? _3919 : _3907;
    assign _3925 = _3913 ? _3924 : _3920;
    assign _3926 = _1058 ? _3925 : _3907;
    assign _3912 = _1055 & _408;
    assign _3927 = _3912 ? _3919 : _3926;
    assign _184 = _3927;
    always @(posedge _416) begin
        if (_414)
            _3907 <= _5492;
        else
            _3907 <= _184;
    end
    assign _3933 = _3932 ? _3907 : _3919;
    assign _3941 = _3929 ? _3940 : _3933;
    assign _3942 = _1058 ? _3941 : _3919;
    assign _3928 = _1055 & _408;
    assign _3943 = _3928 ? _3939 : _3942;
    assign _185 = _3943;
    always @(posedge _416) begin
        if (_414)
            _3919 <= _5492;
        else
            _3919 <= _185;
    end
    assign _3956 = _3955 ? _3919 : _3939;
    assign _3952 = _3948 ? _3951 : _3939;
    assign _3957 = _3945 ? _3956 : _3952;
    assign _3958 = _1058 ? _3957 : _3939;
    assign _3944 = _1055 & _408;
    assign _3959 = _3944 ? _3951 : _3958;
    assign _186 = _3959;
    always @(posedge _416) begin
        if (_414)
            _3939 <= _5492;
        else
            _3939 <= _186;
    end
    assign _3965 = _3964 ? _3939 : _3951;
    assign _3973 = _3961 ? _3972 : _3965;
    assign _3974 = _1058 ? _3973 : _3951;
    assign _3960 = _1055 & _408;
    assign _3975 = _3960 ? _3971 : _3974;
    assign _187 = _3975;
    always @(posedge _416) begin
        if (_414)
            _3951 <= _5492;
        else
            _3951 <= _187;
    end
    assign _3988 = _3987 ? _3951 : _3971;
    assign _3984 = _3980 ? _3983 : _3971;
    assign _3989 = _3977 ? _3988 : _3984;
    assign _3990 = _1058 ? _3989 : _3971;
    assign _3976 = _1055 & _408;
    assign _3991 = _3976 ? _3983 : _3990;
    assign _188 = _3991;
    always @(posedge _416) begin
        if (_414)
            _3971 <= _5492;
        else
            _3971 <= _188;
    end
    assign _3997 = _3996 ? _3971 : _3983;
    assign _4005 = _3993 ? _4004 : _3997;
    assign _4006 = _1058 ? _4005 : _3983;
    assign _3992 = _1055 & _408;
    assign _4007 = _3992 ? _4003 : _4006;
    assign _189 = _4007;
    always @(posedge _416) begin
        if (_414)
            _3983 <= _5492;
        else
            _3983 <= _189;
    end
    assign _4020 = _4019 ? _3983 : _4003;
    assign _4016 = _4012 ? _4015 : _4003;
    assign _4021 = _4009 ? _4020 : _4016;
    assign _4022 = _1058 ? _4021 : _4003;
    assign _4008 = _1055 & _408;
    assign _4023 = _4008 ? _4015 : _4022;
    assign _190 = _4023;
    always @(posedge _416) begin
        if (_414)
            _4003 <= _5492;
        else
            _4003 <= _190;
    end
    assign _4029 = _4028 ? _4003 : _4015;
    assign _4037 = _4025 ? _4036 : _4029;
    assign _4038 = _1058 ? _4037 : _4015;
    assign _4024 = _1055 & _408;
    assign _4039 = _4024 ? _4035 : _4038;
    assign _191 = _4039;
    always @(posedge _416) begin
        if (_414)
            _4015 <= _5492;
        else
            _4015 <= _191;
    end
    assign _4052 = _4051 ? _4015 : _4035;
    assign _4048 = _4044 ? _4047 : _4035;
    assign _4053 = _4041 ? _4052 : _4048;
    assign _4054 = _1058 ? _4053 : _4035;
    assign _4040 = _1055 & _408;
    assign _4055 = _4040 ? _4047 : _4054;
    assign _192 = _4055;
    always @(posedge _416) begin
        if (_414)
            _4035 <= _5492;
        else
            _4035 <= _192;
    end
    assign _4061 = _4060 ? _4035 : _4047;
    assign _4069 = _4057 ? _4068 : _4061;
    assign _4070 = _1058 ? _4069 : _4047;
    assign _4056 = _1055 & _408;
    assign _4071 = _4056 ? _4067 : _4070;
    assign _193 = _4071;
    always @(posedge _416) begin
        if (_414)
            _4047 <= _5492;
        else
            _4047 <= _193;
    end
    assign _4084 = _4083 ? _4047 : _4067;
    assign _4080 = _4076 ? _4079 : _4067;
    assign _4085 = _4073 ? _4084 : _4080;
    assign _4086 = _1058 ? _4085 : _4067;
    assign _4072 = _1055 & _408;
    assign _4087 = _4072 ? _4079 : _4086;
    assign _194 = _4087;
    always @(posedge _416) begin
        if (_414)
            _4067 <= _5492;
        else
            _4067 <= _194;
    end
    assign _4093 = _4092 ? _4067 : _4079;
    assign _4101 = _4089 ? _4100 : _4093;
    assign _4102 = _1058 ? _4101 : _4079;
    assign _4088 = _1055 & _408;
    assign _4103 = _4088 ? _4099 : _4102;
    assign _195 = _4103;
    always @(posedge _416) begin
        if (_414)
            _4079 <= _5492;
        else
            _4079 <= _195;
    end
    assign _4116 = _4115 ? _4079 : _4099;
    assign _4112 = _4108 ? _4111 : _4099;
    assign _4117 = _4105 ? _4116 : _4112;
    assign _4118 = _1058 ? _4117 : _4099;
    assign _4104 = _1055 & _408;
    assign _4119 = _4104 ? _4111 : _4118;
    assign _196 = _4119;
    always @(posedge _416) begin
        if (_414)
            _4099 <= _5492;
        else
            _4099 <= _196;
    end
    assign _4125 = _4124 ? _4099 : _4111;
    assign _4133 = _4121 ? _4132 : _4125;
    assign _4134 = _1058 ? _4133 : _4111;
    assign _4120 = _1055 & _408;
    assign _4135 = _4120 ? _4131 : _4134;
    assign _197 = _4135;
    always @(posedge _416) begin
        if (_414)
            _4111 <= _5492;
        else
            _4111 <= _197;
    end
    assign _4148 = _4147 ? _4111 : _4131;
    assign _4144 = _4140 ? _4143 : _4131;
    assign _4149 = _4137 ? _4148 : _4144;
    assign _4150 = _1058 ? _4149 : _4131;
    assign _4136 = _1055 & _408;
    assign _4151 = _4136 ? _4143 : _4150;
    assign _198 = _4151;
    always @(posedge _416) begin
        if (_414)
            _4131 <= _5492;
        else
            _4131 <= _198;
    end
    assign _4157 = _4156 ? _4131 : _4143;
    assign _4165 = _4153 ? _4164 : _4157;
    assign _4166 = _1058 ? _4165 : _4143;
    assign _4152 = _1055 & _408;
    assign _4167 = _4152 ? _4163 : _4166;
    assign _199 = _4167;
    always @(posedge _416) begin
        if (_414)
            _4143 <= _5492;
        else
            _4143 <= _199;
    end
    assign _4180 = _4179 ? _4143 : _4163;
    assign _4176 = _4172 ? _4175 : _4163;
    assign _4181 = _4169 ? _4180 : _4176;
    assign _4182 = _1058 ? _4181 : _4163;
    assign _4168 = _1055 & _408;
    assign _4183 = _4168 ? _4175 : _4182;
    assign _200 = _4183;
    always @(posedge _416) begin
        if (_414)
            _4163 <= _5492;
        else
            _4163 <= _200;
    end
    assign _4189 = _4188 ? _4163 : _4175;
    assign _4197 = _4185 ? _4196 : _4189;
    assign _4198 = _1058 ? _4197 : _4175;
    assign _4184 = _1055 & _408;
    assign _4199 = _4184 ? _4195 : _4198;
    assign _201 = _4199;
    always @(posedge _416) begin
        if (_414)
            _4175 <= _5492;
        else
            _4175 <= _201;
    end
    assign _4212 = _4211 ? _4175 : _4195;
    assign _4208 = _4204 ? _4207 : _4195;
    assign _4213 = _4201 ? _4212 : _4208;
    assign _4214 = _1058 ? _4213 : _4195;
    assign _4200 = _1055 & _408;
    assign _4215 = _4200 ? _4207 : _4214;
    assign _202 = _4215;
    always @(posedge _416) begin
        if (_414)
            _4195 <= _5492;
        else
            _4195 <= _202;
    end
    assign _4221 = _4220 ? _4195 : _4207;
    assign _4229 = _4217 ? _4228 : _4221;
    assign _4230 = _1058 ? _4229 : _4207;
    assign _4216 = _1055 & _408;
    assign _4231 = _4216 ? _4227 : _4230;
    assign _203 = _4231;
    always @(posedge _416) begin
        if (_414)
            _4207 <= _5492;
        else
            _4207 <= _203;
    end
    assign _4244 = _4243 ? _4207 : _4227;
    assign _4240 = _4236 ? _4239 : _4227;
    assign _4245 = _4233 ? _4244 : _4240;
    assign _4246 = _1058 ? _4245 : _4227;
    assign _4232 = _1055 & _408;
    assign _4247 = _4232 ? _4239 : _4246;
    assign _204 = _4247;
    always @(posedge _416) begin
        if (_414)
            _4227 <= _5492;
        else
            _4227 <= _204;
    end
    assign _5439 = { gnd,
                     _449 };
    assign _4242 = { gnd,
                     _452 };
    assign _4223 = { gnd,
                     _452 };
    assign _4222 = { gnd,
                     _455 };
    assign _4224 = _4222 < _4223;
    assign _5432 = _4224 ? _452 : _455;
    assign _4219 = { gnd,
                     _455 };
    assign _4210 = { gnd,
                     _458 };
    assign _4191 = { gnd,
                     _458 };
    assign _4190 = { gnd,
                     _461 };
    assign _4192 = _4190 < _4191;
    assign _5420 = _4192 ? _458 : _461;
    assign _4187 = { gnd,
                     _461 };
    assign _4178 = { gnd,
                     _464 };
    assign _4159 = { gnd,
                     _464 };
    assign _4158 = { gnd,
                     _467 };
    assign _4160 = _4158 < _4159;
    assign _5408 = _4160 ? _464 : _467;
    assign _4155 = { gnd,
                     _467 };
    assign _4146 = { gnd,
                     _470 };
    assign _4127 = { gnd,
                     _470 };
    assign _4126 = { gnd,
                     _473 };
    assign _4128 = _4126 < _4127;
    assign _5396 = _4128 ? _470 : _473;
    assign _4123 = { gnd,
                     _473 };
    assign _4114 = { gnd,
                     _476 };
    assign _4095 = { gnd,
                     _476 };
    assign _4094 = { gnd,
                     _479 };
    assign _4096 = _4094 < _4095;
    assign _5384 = _4096 ? _476 : _479;
    assign _4091 = { gnd,
                     _479 };
    assign _4082 = { gnd,
                     _482 };
    assign _4063 = { gnd,
                     _482 };
    assign _4062 = { gnd,
                     _485 };
    assign _4064 = _4062 < _4063;
    assign _5372 = _4064 ? _482 : _485;
    assign _4059 = { gnd,
                     _485 };
    assign _4050 = { gnd,
                     _488 };
    assign _4031 = { gnd,
                     _488 };
    assign _4030 = { gnd,
                     _491 };
    assign _4032 = _4030 < _4031;
    assign _5360 = _4032 ? _488 : _491;
    assign _4027 = { gnd,
                     _491 };
    assign _4018 = { gnd,
                     _494 };
    assign _3999 = { gnd,
                     _494 };
    assign _3998 = { gnd,
                     _497 };
    assign _4000 = _3998 < _3999;
    assign _5348 = _4000 ? _494 : _497;
    assign _3995 = { gnd,
                     _497 };
    assign _3986 = { gnd,
                     _500 };
    assign _3967 = { gnd,
                     _500 };
    assign _3966 = { gnd,
                     _503 };
    assign _3968 = _3966 < _3967;
    assign _5336 = _3968 ? _500 : _503;
    assign _3963 = { gnd,
                     _503 };
    assign _3954 = { gnd,
                     _506 };
    assign _3935 = { gnd,
                     _506 };
    assign _3934 = { gnd,
                     _509 };
    assign _3936 = _3934 < _3935;
    assign _5324 = _3936 ? _506 : _509;
    assign _3931 = { gnd,
                     _509 };
    assign _3922 = { gnd,
                     _512 };
    assign _3903 = { gnd,
                     _512 };
    assign _3902 = { gnd,
                     _515 };
    assign _3904 = _3902 < _3903;
    assign _5312 = _3904 ? _512 : _515;
    assign _3899 = { gnd,
                     _515 };
    assign _3890 = { gnd,
                     _518 };
    assign _3871 = { gnd,
                     _518 };
    assign _3870 = { gnd,
                     _521 };
    assign _3872 = _3870 < _3871;
    assign _5300 = _3872 ? _518 : _521;
    assign _3867 = { gnd,
                     _521 };
    assign _3858 = { gnd,
                     _524 };
    assign _3839 = { gnd,
                     _524 };
    assign _3838 = { gnd,
                     _527 };
    assign _3840 = _3838 < _3839;
    assign _5288 = _3840 ? _524 : _527;
    assign _3835 = { gnd,
                     _527 };
    assign _3826 = { gnd,
                     _530 };
    assign _3807 = { gnd,
                     _530 };
    assign _3806 = { gnd,
                     _533 };
    assign _3808 = _3806 < _3807;
    assign _5276 = _3808 ? _530 : _533;
    assign _3803 = { gnd,
                     _533 };
    assign _3794 = { gnd,
                     _536 };
    assign _3775 = { gnd,
                     _536 };
    assign _3774 = { gnd,
                     _539 };
    assign _3776 = _3774 < _3775;
    assign _5264 = _3776 ? _536 : _539;
    assign _3771 = { gnd,
                     _539 };
    assign _3762 = { gnd,
                     _542 };
    assign _3743 = { gnd,
                     _542 };
    assign _3742 = { gnd,
                     _545 };
    assign _3744 = _3742 < _3743;
    assign _5252 = _3744 ? _542 : _545;
    assign _3739 = { gnd,
                     _545 };
    assign _3730 = { gnd,
                     _548 };
    assign _3711 = { gnd,
                     _548 };
    assign _3710 = { gnd,
                     _551 };
    assign _3712 = _3710 < _3711;
    assign _5240 = _3712 ? _548 : _551;
    assign _3707 = { gnd,
                     _551 };
    assign _3698 = { gnd,
                     _554 };
    assign _3679 = { gnd,
                     _554 };
    assign _3678 = { gnd,
                     _557 };
    assign _3680 = _3678 < _3679;
    assign _5228 = _3680 ? _554 : _557;
    assign _3675 = { gnd,
                     _557 };
    assign _3666 = { gnd,
                     _560 };
    assign _3647 = { gnd,
                     _560 };
    assign _3646 = { gnd,
                     _563 };
    assign _3648 = _3646 < _3647;
    assign _5216 = _3648 ? _560 : _563;
    assign _3643 = { gnd,
                     _563 };
    assign _3634 = { gnd,
                     _566 };
    assign _3615 = { gnd,
                     _566 };
    assign _3614 = { gnd,
                     _569 };
    assign _3616 = _3614 < _3615;
    assign _5204 = _3616 ? _566 : _569;
    assign _3611 = { gnd,
                     _569 };
    assign _3602 = { gnd,
                     _572 };
    assign _3583 = { gnd,
                     _572 };
    assign _3582 = { gnd,
                     _575 };
    assign _3584 = _3582 < _3583;
    assign _5192 = _3584 ? _572 : _575;
    assign _3579 = { gnd,
                     _575 };
    assign _3570 = { gnd,
                     _578 };
    assign _3551 = { gnd,
                     _578 };
    assign _3550 = { gnd,
                     _581 };
    assign _3552 = _3550 < _3551;
    assign _5180 = _3552 ? _578 : _581;
    assign _3547 = { gnd,
                     _581 };
    assign _3538 = { gnd,
                     _584 };
    assign _3519 = { gnd,
                     _584 };
    assign _3518 = { gnd,
                     _587 };
    assign _3520 = _3518 < _3519;
    assign _5168 = _3520 ? _584 : _587;
    assign _3515 = { gnd,
                     _587 };
    assign _3506 = { gnd,
                     _590 };
    assign _3487 = { gnd,
                     _590 };
    assign _3486 = { gnd,
                     _593 };
    assign _3488 = _3486 < _3487;
    assign _5156 = _3488 ? _590 : _593;
    assign _3483 = { gnd,
                     _593 };
    assign _3474 = { gnd,
                     _596 };
    assign _3455 = { gnd,
                     _596 };
    assign _3454 = { gnd,
                     _599 };
    assign _3456 = _3454 < _3455;
    assign _5144 = _3456 ? _596 : _599;
    assign _3451 = { gnd,
                     _599 };
    assign _3442 = { gnd,
                     _602 };
    assign _3423 = { gnd,
                     _602 };
    assign _3422 = { gnd,
                     _605 };
    assign _3424 = _3422 < _3423;
    assign _5132 = _3424 ? _602 : _605;
    assign _3419 = { gnd,
                     _605 };
    assign _3410 = { gnd,
                     _608 };
    assign _3391 = { gnd,
                     _608 };
    assign _3390 = { gnd,
                     _611 };
    assign _3392 = _3390 < _3391;
    assign _5120 = _3392 ? _608 : _611;
    assign _3387 = { gnd,
                     _611 };
    assign _3378 = { gnd,
                     _614 };
    assign _3359 = { gnd,
                     _614 };
    assign _3358 = { gnd,
                     _617 };
    assign _3360 = _3358 < _3359;
    assign _5108 = _3360 ? _614 : _617;
    assign _3355 = { gnd,
                     _617 };
    assign _3346 = { gnd,
                     _620 };
    assign _3327 = { gnd,
                     _620 };
    assign _3326 = { gnd,
                     _623 };
    assign _3328 = _3326 < _3327;
    assign _5096 = _3328 ? _620 : _623;
    assign _3323 = { gnd,
                     _623 };
    assign _3314 = { gnd,
                     _626 };
    assign _3295 = { gnd,
                     _626 };
    assign _3294 = { gnd,
                     _629 };
    assign _3296 = _3294 < _3295;
    assign _5084 = _3296 ? _626 : _629;
    assign _3291 = { gnd,
                     _629 };
    assign _3282 = { gnd,
                     _632 };
    assign _3263 = { gnd,
                     _632 };
    assign _3262 = { gnd,
                     _635 };
    assign _3264 = _3262 < _3263;
    assign _5072 = _3264 ? _632 : _635;
    assign _3259 = { gnd,
                     _635 };
    assign _3250 = { gnd,
                     _638 };
    assign _3231 = { gnd,
                     _638 };
    assign _3230 = { gnd,
                     _641 };
    assign _3232 = _3230 < _3231;
    assign _5060 = _3232 ? _638 : _641;
    assign _3227 = { gnd,
                     _641 };
    assign _3218 = { gnd,
                     _644 };
    assign _3199 = { gnd,
                     _644 };
    assign _3198 = { gnd,
                     _647 };
    assign _3200 = _3198 < _3199;
    assign _5048 = _3200 ? _644 : _647;
    assign _3195 = { gnd,
                     _647 };
    assign _3186 = { gnd,
                     _650 };
    assign _3167 = { gnd,
                     _650 };
    assign _3166 = { gnd,
                     _653 };
    assign _3168 = _3166 < _3167;
    assign _5036 = _3168 ? _650 : _653;
    assign _3163 = { gnd,
                     _653 };
    assign _3154 = { gnd,
                     _656 };
    assign _3135 = { gnd,
                     _656 };
    assign _3134 = { gnd,
                     _659 };
    assign _3136 = _3134 < _3135;
    assign _5024 = _3136 ? _656 : _659;
    assign _3131 = { gnd,
                     _659 };
    assign _3122 = { gnd,
                     _662 };
    assign _3103 = { gnd,
                     _662 };
    assign _3102 = { gnd,
                     _665 };
    assign _3104 = _3102 < _3103;
    assign _5012 = _3104 ? _662 : _665;
    assign _3099 = { gnd,
                     _665 };
    assign _3090 = { gnd,
                     _668 };
    assign _3071 = { gnd,
                     _668 };
    assign _3070 = { gnd,
                     _671 };
    assign _3072 = _3070 < _3071;
    assign _5000 = _3072 ? _668 : _671;
    assign _3067 = { gnd,
                     _671 };
    assign _3058 = { gnd,
                     _674 };
    assign _3039 = { gnd,
                     _674 };
    assign _3038 = { gnd,
                     _677 };
    assign _3040 = _3038 < _3039;
    assign _4988 = _3040 ? _674 : _677;
    assign _3035 = { gnd,
                     _677 };
    assign _3026 = { gnd,
                     _680 };
    assign _3007 = { gnd,
                     _680 };
    assign _3006 = { gnd,
                     _683 };
    assign _3008 = _3006 < _3007;
    assign _4976 = _3008 ? _680 : _683;
    assign _3003 = { gnd,
                     _683 };
    assign _2994 = { gnd,
                     _686 };
    assign _2975 = { gnd,
                     _686 };
    assign _2974 = { gnd,
                     _689 };
    assign _2976 = _2974 < _2975;
    assign _4964 = _2976 ? _686 : _689;
    assign _2971 = { gnd,
                     _689 };
    assign _2962 = { gnd,
                     _692 };
    assign _2943 = { gnd,
                     _692 };
    assign _2942 = { gnd,
                     _695 };
    assign _2944 = _2942 < _2943;
    assign _4952 = _2944 ? _692 : _695;
    assign _2939 = { gnd,
                     _695 };
    assign _2930 = { gnd,
                     _698 };
    assign _2911 = { gnd,
                     _698 };
    assign _2910 = { gnd,
                     _701 };
    assign _2912 = _2910 < _2911;
    assign _4940 = _2912 ? _698 : _701;
    assign _2907 = { gnd,
                     _701 };
    assign _2898 = { gnd,
                     _704 };
    assign _2879 = { gnd,
                     _704 };
    assign _2878 = { gnd,
                     _707 };
    assign _2880 = _2878 < _2879;
    assign _4928 = _2880 ? _704 : _707;
    assign _2875 = { gnd,
                     _707 };
    assign _2866 = { gnd,
                     _710 };
    assign _2847 = { gnd,
                     _710 };
    assign _2846 = { gnd,
                     _713 };
    assign _2848 = _2846 < _2847;
    assign _4916 = _2848 ? _710 : _713;
    assign _2843 = { gnd,
                     _713 };
    assign _2834 = { gnd,
                     _716 };
    assign _2815 = { gnd,
                     _716 };
    assign _2814 = { gnd,
                     _719 };
    assign _2816 = _2814 < _2815;
    assign _4904 = _2816 ? _716 : _719;
    assign _2811 = { gnd,
                     _719 };
    assign _2802 = { gnd,
                     _722 };
    assign _2783 = { gnd,
                     _722 };
    assign _2782 = { gnd,
                     _725 };
    assign _2784 = _2782 < _2783;
    assign _4892 = _2784 ? _722 : _725;
    assign _2779 = { gnd,
                     _725 };
    assign _2770 = { gnd,
                     _728 };
    assign _2751 = { gnd,
                     _728 };
    assign _2750 = { gnd,
                     _731 };
    assign _2752 = _2750 < _2751;
    assign _4880 = _2752 ? _728 : _731;
    assign _2747 = { gnd,
                     _731 };
    assign _2738 = { gnd,
                     _734 };
    assign _2719 = { gnd,
                     _734 };
    assign _2718 = { gnd,
                     _737 };
    assign _2720 = _2718 < _2719;
    assign _4868 = _2720 ? _734 : _737;
    assign _2715 = { gnd,
                     _737 };
    assign _2706 = { gnd,
                     _740 };
    assign _2687 = { gnd,
                     _740 };
    assign _2686 = { gnd,
                     _743 };
    assign _2688 = _2686 < _2687;
    assign _4856 = _2688 ? _740 : _743;
    assign _2683 = { gnd,
                     _743 };
    assign _2674 = { gnd,
                     _746 };
    assign _2655 = { gnd,
                     _746 };
    assign _2654 = { gnd,
                     _749 };
    assign _2656 = _2654 < _2655;
    assign _4844 = _2656 ? _746 : _749;
    assign _2651 = { gnd,
                     _749 };
    assign _2642 = { gnd,
                     _752 };
    assign _2623 = { gnd,
                     _752 };
    assign _2622 = { gnd,
                     _755 };
    assign _2624 = _2622 < _2623;
    assign _4832 = _2624 ? _752 : _755;
    assign _2619 = { gnd,
                     _755 };
    assign _2610 = { gnd,
                     _758 };
    assign _2591 = { gnd,
                     _758 };
    assign _2590 = { gnd,
                     _761 };
    assign _2592 = _2590 < _2591;
    assign _4820 = _2592 ? _758 : _761;
    assign _2587 = { gnd,
                     _761 };
    assign _2578 = { gnd,
                     _764 };
    assign _2559 = { gnd,
                     _764 };
    assign _2558 = { gnd,
                     _767 };
    assign _2560 = _2558 < _2559;
    assign _4808 = _2560 ? _764 : _767;
    assign _2555 = { gnd,
                     _767 };
    assign _2546 = { gnd,
                     _770 };
    assign _2527 = { gnd,
                     _770 };
    assign _2526 = { gnd,
                     _773 };
    assign _2528 = _2526 < _2527;
    assign _4796 = _2528 ? _770 : _773;
    assign _2523 = { gnd,
                     _773 };
    assign _2514 = { gnd,
                     _776 };
    assign _2495 = { gnd,
                     _776 };
    assign _2494 = { gnd,
                     _779 };
    assign _2496 = _2494 < _2495;
    assign _4784 = _2496 ? _776 : _779;
    assign _2491 = { gnd,
                     _779 };
    assign _2482 = { gnd,
                     _782 };
    assign _2463 = { gnd,
                     _782 };
    assign _2462 = { gnd,
                     _785 };
    assign _2464 = _2462 < _2463;
    assign _4772 = _2464 ? _782 : _785;
    assign _2459 = { gnd,
                     _785 };
    assign _2450 = { gnd,
                     _788 };
    assign _2431 = { gnd,
                     _788 };
    assign _2430 = { gnd,
                     _791 };
    assign _2432 = _2430 < _2431;
    assign _4760 = _2432 ? _788 : _791;
    assign _2427 = { gnd,
                     _791 };
    assign _2418 = { gnd,
                     _794 };
    assign _2399 = { gnd,
                     _794 };
    assign _2398 = { gnd,
                     _797 };
    assign _2400 = _2398 < _2399;
    assign _4748 = _2400 ? _794 : _797;
    assign _2395 = { gnd,
                     _797 };
    assign _2386 = { gnd,
                     _800 };
    assign _2367 = { gnd,
                     _800 };
    assign _2366 = { gnd,
                     _803 };
    assign _2368 = _2366 < _2367;
    assign _4736 = _2368 ? _800 : _803;
    assign _2363 = { gnd,
                     _803 };
    assign _2354 = { gnd,
                     _806 };
    assign _2335 = { gnd,
                     _806 };
    assign _2334 = { gnd,
                     _809 };
    assign _2336 = _2334 < _2335;
    assign _4724 = _2336 ? _806 : _809;
    assign _2331 = { gnd,
                     _809 };
    assign _2322 = { gnd,
                     _812 };
    assign _2303 = { gnd,
                     _812 };
    assign _2302 = { gnd,
                     _815 };
    assign _2304 = _2302 < _2303;
    assign _4712 = _2304 ? _812 : _815;
    assign _2299 = { gnd,
                     _815 };
    assign _2290 = { gnd,
                     _818 };
    assign _2271 = { gnd,
                     _818 };
    assign _2270 = { gnd,
                     _821 };
    assign _2272 = _2270 < _2271;
    assign _4700 = _2272 ? _818 : _821;
    assign _2267 = { gnd,
                     _821 };
    assign _2258 = { gnd,
                     _824 };
    assign _2239 = { gnd,
                     _824 };
    assign _2238 = { gnd,
                     _827 };
    assign _2240 = _2238 < _2239;
    assign _4688 = _2240 ? _824 : _827;
    assign _2235 = { gnd,
                     _827 };
    assign _2226 = { gnd,
                     _830 };
    assign _2207 = { gnd,
                     _830 };
    assign _2206 = { gnd,
                     _833 };
    assign _2208 = _2206 < _2207;
    assign _4676 = _2208 ? _830 : _833;
    assign _2203 = { gnd,
                     _833 };
    assign _2194 = { gnd,
                     _836 };
    assign _2175 = { gnd,
                     _836 };
    assign _2174 = { gnd,
                     _839 };
    assign _2176 = _2174 < _2175;
    assign _4664 = _2176 ? _836 : _839;
    assign _2171 = { gnd,
                     _839 };
    assign _2162 = { gnd,
                     _842 };
    assign _2143 = { gnd,
                     _842 };
    assign _2142 = { gnd,
                     _845 };
    assign _2144 = _2142 < _2143;
    assign _4652 = _2144 ? _842 : _845;
    assign _2139 = { gnd,
                     _845 };
    assign _2130 = { gnd,
                     _848 };
    assign _2111 = { gnd,
                     _848 };
    assign _2110 = { gnd,
                     _851 };
    assign _2112 = _2110 < _2111;
    assign _4640 = _2112 ? _848 : _851;
    assign _2107 = { gnd,
                     _851 };
    assign _2098 = { gnd,
                     _854 };
    assign _2079 = { gnd,
                     _854 };
    assign _2078 = { gnd,
                     _857 };
    assign _2080 = _2078 < _2079;
    assign _4628 = _2080 ? _854 : _857;
    assign _2075 = { gnd,
                     _857 };
    assign _2066 = { gnd,
                     _860 };
    assign _2047 = { gnd,
                     _860 };
    assign _2046 = { gnd,
                     _863 };
    assign _2048 = _2046 < _2047;
    assign _4616 = _2048 ? _860 : _863;
    assign _2043 = { gnd,
                     _863 };
    assign _2034 = { gnd,
                     _866 };
    assign _2015 = { gnd,
                     _866 };
    assign _2014 = { gnd,
                     _869 };
    assign _2016 = _2014 < _2015;
    assign _4604 = _2016 ? _866 : _869;
    assign _2011 = { gnd,
                     _869 };
    assign _2002 = { gnd,
                     _872 };
    assign _1983 = { gnd,
                     _872 };
    assign _1982 = { gnd,
                     _875 };
    assign _1984 = _1982 < _1983;
    assign _4592 = _1984 ? _872 : _875;
    assign _1979 = { gnd,
                     _875 };
    assign _1970 = { gnd,
                     _878 };
    assign _1951 = { gnd,
                     _878 };
    assign _1950 = { gnd,
                     _881 };
    assign _1952 = _1950 < _1951;
    assign _4580 = _1952 ? _878 : _881;
    assign _1947 = { gnd,
                     _881 };
    assign _1938 = { gnd,
                     _884 };
    assign _1919 = { gnd,
                     _884 };
    assign _1918 = { gnd,
                     _887 };
    assign _1920 = _1918 < _1919;
    assign _4568 = _1920 ? _884 : _887;
    assign _1915 = { gnd,
                     _887 };
    assign _1906 = { gnd,
                     _890 };
    assign _1887 = { gnd,
                     _890 };
    assign _1886 = { gnd,
                     _893 };
    assign _1888 = _1886 < _1887;
    assign _4556 = _1888 ? _890 : _893;
    assign _1883 = { gnd,
                     _893 };
    assign _1874 = { gnd,
                     _896 };
    assign _1855 = { gnd,
                     _896 };
    assign _1854 = { gnd,
                     _899 };
    assign _1856 = _1854 < _1855;
    assign _4544 = _1856 ? _896 : _899;
    assign _1851 = { gnd,
                     _899 };
    assign _1842 = { gnd,
                     _902 };
    assign _1823 = { gnd,
                     _902 };
    assign _1822 = { gnd,
                     _905 };
    assign _1824 = _1822 < _1823;
    assign _4532 = _1824 ? _902 : _905;
    assign _1819 = { gnd,
                     _905 };
    assign _1810 = { gnd,
                     _908 };
    assign _1791 = { gnd,
                     _908 };
    assign _1790 = { gnd,
                     _911 };
    assign _1792 = _1790 < _1791;
    assign _4520 = _1792 ? _908 : _911;
    assign _1787 = { gnd,
                     _911 };
    assign _1778 = { gnd,
                     _914 };
    assign _1759 = { gnd,
                     _914 };
    assign _1758 = { gnd,
                     _917 };
    assign _1760 = _1758 < _1759;
    assign _4508 = _1760 ? _914 : _917;
    assign _1755 = { gnd,
                     _917 };
    assign _1746 = { gnd,
                     _920 };
    assign _1727 = { gnd,
                     _920 };
    assign _1726 = { gnd,
                     _923 };
    assign _1728 = _1726 < _1727;
    assign _4496 = _1728 ? _920 : _923;
    assign _1723 = { gnd,
                     _923 };
    assign _1714 = { gnd,
                     _926 };
    assign _1695 = { gnd,
                     _926 };
    assign _1694 = { gnd,
                     _929 };
    assign _1696 = _1694 < _1695;
    assign _4484 = _1696 ? _926 : _929;
    assign _1691 = { gnd,
                     _929 };
    assign _1682 = { gnd,
                     _932 };
    assign _1663 = { gnd,
                     _932 };
    assign _1662 = { gnd,
                     _935 };
    assign _1664 = _1662 < _1663;
    assign _4472 = _1664 ? _932 : _935;
    assign _1659 = { gnd,
                     _935 };
    assign _1650 = { gnd,
                     _938 };
    assign _1631 = { gnd,
                     _938 };
    assign _1630 = { gnd,
                     _941 };
    assign _1632 = _1630 < _1631;
    assign _4460 = _1632 ? _938 : _941;
    assign _1627 = { gnd,
                     _941 };
    assign _1618 = { gnd,
                     _944 };
    assign _1599 = { gnd,
                     _944 };
    assign _1598 = { gnd,
                     _947 };
    assign _1600 = _1598 < _1599;
    assign _4448 = _1600 ? _944 : _947;
    assign _1595 = { gnd,
                     _947 };
    assign _1586 = { gnd,
                     _950 };
    assign _1567 = { gnd,
                     _950 };
    assign _1566 = { gnd,
                     _953 };
    assign _1568 = _1566 < _1567;
    assign _4436 = _1568 ? _950 : _953;
    assign _1563 = { gnd,
                     _953 };
    assign _1554 = { gnd,
                     _956 };
    assign _1535 = { gnd,
                     _956 };
    assign _1534 = { gnd,
                     _959 };
    assign _1536 = _1534 < _1535;
    assign _4424 = _1536 ? _956 : _959;
    assign _1531 = { gnd,
                     _959 };
    assign _1522 = { gnd,
                     _962 };
    assign _1503 = { gnd,
                     _962 };
    assign _1502 = { gnd,
                     _965 };
    assign _1504 = _1502 < _1503;
    assign _4412 = _1504 ? _962 : _965;
    assign _1499 = { gnd,
                     _965 };
    assign _1490 = { gnd,
                     _968 };
    assign _1471 = { gnd,
                     _968 };
    assign _1470 = { gnd,
                     _971 };
    assign _1472 = _1470 < _1471;
    assign _4400 = _1472 ? _968 : _971;
    assign _1467 = { gnd,
                     _971 };
    assign _1458 = { gnd,
                     _974 };
    assign _1439 = { gnd,
                     _974 };
    assign _1438 = { gnd,
                     _977 };
    assign _1440 = _1438 < _1439;
    assign _4388 = _1440 ? _974 : _977;
    assign _1435 = { gnd,
                     _977 };
    assign _1426 = { gnd,
                     _980 };
    assign _1407 = { gnd,
                     _980 };
    assign _1406 = { gnd,
                     _983 };
    assign _1408 = _1406 < _1407;
    assign _4376 = _1408 ? _980 : _983;
    assign _1403 = { gnd,
                     _983 };
    assign _1394 = { gnd,
                     _986 };
    assign _1375 = { gnd,
                     _986 };
    assign _1374 = { gnd,
                     _989 };
    assign _1376 = _1374 < _1375;
    assign _4364 = _1376 ? _986 : _989;
    assign _1371 = { gnd,
                     _989 };
    assign _1362 = { gnd,
                     _992 };
    assign _1343 = { gnd,
                     _992 };
    assign _1342 = { gnd,
                     _995 };
    assign _1344 = _1342 < _1343;
    assign _4352 = _1344 ? _992 : _995;
    assign _1339 = { gnd,
                     _995 };
    assign _1330 = { gnd,
                     _998 };
    assign _1311 = { gnd,
                     _998 };
    assign _1310 = { gnd,
                     _1001 };
    assign _1312 = _1310 < _1311;
    assign _4340 = _1312 ? _998 : _1001;
    assign _1307 = { gnd,
                     _1001 };
    assign _1298 = { gnd,
                     _1004 };
    assign _1279 = { gnd,
                     _1004 };
    assign _1278 = { gnd,
                     _1007 };
    assign _1280 = _1278 < _1279;
    assign _4328 = _1280 ? _1004 : _1007;
    assign _1275 = { gnd,
                     _1007 };
    assign _1266 = { gnd,
                     _1010 };
    assign _1247 = { gnd,
                     _1010 };
    assign _1246 = { gnd,
                     _1013 };
    assign _1248 = _1246 < _1247;
    assign _4316 = _1248 ? _1010 : _1013;
    assign _1243 = { gnd,
                     _1013 };
    assign _1234 = { gnd,
                     _1016 };
    assign _1215 = { gnd,
                     _1016 };
    assign _1214 = { gnd,
                     _1019 };
    assign _1216 = _1214 < _1215;
    assign _4304 = _1216 ? _1016 : _1019;
    assign _1211 = { gnd,
                     _1019 };
    assign _1202 = { gnd,
                     _1022 };
    assign _1183 = { gnd,
                     _1022 };
    assign _1182 = { gnd,
                     _1025 };
    assign _1184 = _1182 < _1183;
    assign _4292 = _1184 ? _1022 : _1025;
    assign _1179 = { gnd,
                     _1025 };
    assign _1170 = { gnd,
                     _1028 };
    assign _1151 = { gnd,
                     _1028 };
    assign _1150 = { gnd,
                     _1031 };
    assign _1152 = _1150 < _1151;
    assign _4280 = _1152 ? _1028 : _1031;
    assign _1147 = { gnd,
                     _1031 };
    assign _1138 = { gnd,
                     _1034 };
    assign _1119 = { gnd,
                     _1034 };
    assign _1118 = { gnd,
                     _1037 };
    assign _1120 = _1118 < _1119;
    assign _4268 = _1120 ? _1034 : _1037;
    assign _1115 = { gnd,
                     _1037 };
    assign _1106 = { gnd,
                     _1040 };
    assign _1087 = { gnd,
                     _1040 };
    assign _1086 = { gnd,
                     _1043 };
    assign _1088 = _1086 < _1087;
    assign _4256 = _1088 ? _1040 : _1043;
    assign _1083 = { gnd,
                     _1043 };
    assign _1074 = { gnd,
                     _1046 };
    assign _1073 = { gnd,
                     _1046 };
    assign _1075 = _1073 < _1074;
    assign _4250 = _1075 ? _1046 : _1046;
    assign _1067 = { gnd,
                     _1043 };
    assign _1066 = { gnd,
                     _1046 };
    assign _1068 = _1066 < _1067;
    assign _4249 = _1068 ? _1043 : _1046;
    assign _1065 = _1064[0:0];
    assign _4251 = _1065 ? _4250 : _4249;
    assign _4252 = _1058 ? _4251 : _1046;
    assign _4248 = _1055 & _408;
    assign _4253 = _4248 ? _1043 : _4252;
    assign _205 = _4253;
    always @(posedge _416) begin
        if (_414)
            _1046 <= _5492;
        else
            _1046 <= _205;
    end
    assign _1082 = { gnd,
                     _1046 };
    assign _1084 = _1082 < _1083;
    assign _4255 = _1084 ? _1046 : _1043;
    assign _1081 = _1064[0:0];
    assign _4257 = _1081 ? _4256 : _4255;
    assign _4258 = _1058 ? _4257 : _1043;
    assign _4254 = _1055 & _408;
    assign _4259 = _4254 ? _1040 : _4258;
    assign _206 = _4259;
    always @(posedge _416) begin
        if (_414)
            _1043 <= _5492;
        else
            _1043 <= _206;
    end
    assign _1105 = { gnd,
                     _1043 };
    assign _1107 = _1105 < _1106;
    assign _4262 = _1107 ? _1043 : _1040;
    assign _1099 = { gnd,
                     _1037 };
    assign _1098 = { gnd,
                     _1040 };
    assign _1100 = _1098 < _1099;
    assign _4261 = _1100 ? _1037 : _1040;
    assign _1097 = _1064[0:0];
    assign _4263 = _1097 ? _4262 : _4261;
    assign _4264 = _1058 ? _4263 : _1040;
    assign _4260 = _1055 & _408;
    assign _4265 = _4260 ? _1037 : _4264;
    assign _207 = _4265;
    always @(posedge _416) begin
        if (_414)
            _1040 <= _5492;
        else
            _1040 <= _207;
    end
    assign _1114 = { gnd,
                     _1040 };
    assign _1116 = _1114 < _1115;
    assign _4267 = _1116 ? _1040 : _1037;
    assign _1113 = _1064[0:0];
    assign _4269 = _1113 ? _4268 : _4267;
    assign _4270 = _1058 ? _4269 : _1037;
    assign _4266 = _1055 & _408;
    assign _4271 = _4266 ? _1034 : _4270;
    assign _208 = _4271;
    always @(posedge _416) begin
        if (_414)
            _1037 <= _5492;
        else
            _1037 <= _208;
    end
    assign _1137 = { gnd,
                     _1037 };
    assign _1139 = _1137 < _1138;
    assign _4274 = _1139 ? _1037 : _1034;
    assign _1131 = { gnd,
                     _1031 };
    assign _1130 = { gnd,
                     _1034 };
    assign _1132 = _1130 < _1131;
    assign _4273 = _1132 ? _1031 : _1034;
    assign _1129 = _1064[0:0];
    assign _4275 = _1129 ? _4274 : _4273;
    assign _4276 = _1058 ? _4275 : _1034;
    assign _4272 = _1055 & _408;
    assign _4277 = _4272 ? _1031 : _4276;
    assign _209 = _4277;
    always @(posedge _416) begin
        if (_414)
            _1034 <= _5492;
        else
            _1034 <= _209;
    end
    assign _1146 = { gnd,
                     _1034 };
    assign _1148 = _1146 < _1147;
    assign _4279 = _1148 ? _1034 : _1031;
    assign _1145 = _1064[0:0];
    assign _4281 = _1145 ? _4280 : _4279;
    assign _4282 = _1058 ? _4281 : _1031;
    assign _4278 = _1055 & _408;
    assign _4283 = _4278 ? _1028 : _4282;
    assign _210 = _4283;
    always @(posedge _416) begin
        if (_414)
            _1031 <= _5492;
        else
            _1031 <= _210;
    end
    assign _1169 = { gnd,
                     _1031 };
    assign _1171 = _1169 < _1170;
    assign _4286 = _1171 ? _1031 : _1028;
    assign _1163 = { gnd,
                     _1025 };
    assign _1162 = { gnd,
                     _1028 };
    assign _1164 = _1162 < _1163;
    assign _4285 = _1164 ? _1025 : _1028;
    assign _1161 = _1064[0:0];
    assign _4287 = _1161 ? _4286 : _4285;
    assign _4288 = _1058 ? _4287 : _1028;
    assign _4284 = _1055 & _408;
    assign _4289 = _4284 ? _1025 : _4288;
    assign _211 = _4289;
    always @(posedge _416) begin
        if (_414)
            _1028 <= _5492;
        else
            _1028 <= _211;
    end
    assign _1178 = { gnd,
                     _1028 };
    assign _1180 = _1178 < _1179;
    assign _4291 = _1180 ? _1028 : _1025;
    assign _1177 = _1064[0:0];
    assign _4293 = _1177 ? _4292 : _4291;
    assign _4294 = _1058 ? _4293 : _1025;
    assign _4290 = _1055 & _408;
    assign _4295 = _4290 ? _1022 : _4294;
    assign _212 = _4295;
    always @(posedge _416) begin
        if (_414)
            _1025 <= _5492;
        else
            _1025 <= _212;
    end
    assign _1201 = { gnd,
                     _1025 };
    assign _1203 = _1201 < _1202;
    assign _4298 = _1203 ? _1025 : _1022;
    assign _1195 = { gnd,
                     _1019 };
    assign _1194 = { gnd,
                     _1022 };
    assign _1196 = _1194 < _1195;
    assign _4297 = _1196 ? _1019 : _1022;
    assign _1193 = _1064[0:0];
    assign _4299 = _1193 ? _4298 : _4297;
    assign _4300 = _1058 ? _4299 : _1022;
    assign _4296 = _1055 & _408;
    assign _4301 = _4296 ? _1019 : _4300;
    assign _213 = _4301;
    always @(posedge _416) begin
        if (_414)
            _1022 <= _5492;
        else
            _1022 <= _213;
    end
    assign _1210 = { gnd,
                     _1022 };
    assign _1212 = _1210 < _1211;
    assign _4303 = _1212 ? _1022 : _1019;
    assign _1209 = _1064[0:0];
    assign _4305 = _1209 ? _4304 : _4303;
    assign _4306 = _1058 ? _4305 : _1019;
    assign _4302 = _1055 & _408;
    assign _4307 = _4302 ? _1016 : _4306;
    assign _214 = _4307;
    always @(posedge _416) begin
        if (_414)
            _1019 <= _5492;
        else
            _1019 <= _214;
    end
    assign _1233 = { gnd,
                     _1019 };
    assign _1235 = _1233 < _1234;
    assign _4310 = _1235 ? _1019 : _1016;
    assign _1227 = { gnd,
                     _1013 };
    assign _1226 = { gnd,
                     _1016 };
    assign _1228 = _1226 < _1227;
    assign _4309 = _1228 ? _1013 : _1016;
    assign _1225 = _1064[0:0];
    assign _4311 = _1225 ? _4310 : _4309;
    assign _4312 = _1058 ? _4311 : _1016;
    assign _4308 = _1055 & _408;
    assign _4313 = _4308 ? _1013 : _4312;
    assign _215 = _4313;
    always @(posedge _416) begin
        if (_414)
            _1016 <= _5492;
        else
            _1016 <= _215;
    end
    assign _1242 = { gnd,
                     _1016 };
    assign _1244 = _1242 < _1243;
    assign _4315 = _1244 ? _1016 : _1013;
    assign _1241 = _1064[0:0];
    assign _4317 = _1241 ? _4316 : _4315;
    assign _4318 = _1058 ? _4317 : _1013;
    assign _4314 = _1055 & _408;
    assign _4319 = _4314 ? _1010 : _4318;
    assign _216 = _4319;
    always @(posedge _416) begin
        if (_414)
            _1013 <= _5492;
        else
            _1013 <= _216;
    end
    assign _1265 = { gnd,
                     _1013 };
    assign _1267 = _1265 < _1266;
    assign _4322 = _1267 ? _1013 : _1010;
    assign _1259 = { gnd,
                     _1007 };
    assign _1258 = { gnd,
                     _1010 };
    assign _1260 = _1258 < _1259;
    assign _4321 = _1260 ? _1007 : _1010;
    assign _1257 = _1064[0:0];
    assign _4323 = _1257 ? _4322 : _4321;
    assign _4324 = _1058 ? _4323 : _1010;
    assign _4320 = _1055 & _408;
    assign _4325 = _4320 ? _1007 : _4324;
    assign _217 = _4325;
    always @(posedge _416) begin
        if (_414)
            _1010 <= _5492;
        else
            _1010 <= _217;
    end
    assign _1274 = { gnd,
                     _1010 };
    assign _1276 = _1274 < _1275;
    assign _4327 = _1276 ? _1010 : _1007;
    assign _1273 = _1064[0:0];
    assign _4329 = _1273 ? _4328 : _4327;
    assign _4330 = _1058 ? _4329 : _1007;
    assign _4326 = _1055 & _408;
    assign _4331 = _4326 ? _1004 : _4330;
    assign _218 = _4331;
    always @(posedge _416) begin
        if (_414)
            _1007 <= _5492;
        else
            _1007 <= _218;
    end
    assign _1297 = { gnd,
                     _1007 };
    assign _1299 = _1297 < _1298;
    assign _4334 = _1299 ? _1007 : _1004;
    assign _1291 = { gnd,
                     _1001 };
    assign _1290 = { gnd,
                     _1004 };
    assign _1292 = _1290 < _1291;
    assign _4333 = _1292 ? _1001 : _1004;
    assign _1289 = _1064[0:0];
    assign _4335 = _1289 ? _4334 : _4333;
    assign _4336 = _1058 ? _4335 : _1004;
    assign _4332 = _1055 & _408;
    assign _4337 = _4332 ? _1001 : _4336;
    assign _219 = _4337;
    always @(posedge _416) begin
        if (_414)
            _1004 <= _5492;
        else
            _1004 <= _219;
    end
    assign _1306 = { gnd,
                     _1004 };
    assign _1308 = _1306 < _1307;
    assign _4339 = _1308 ? _1004 : _1001;
    assign _1305 = _1064[0:0];
    assign _4341 = _1305 ? _4340 : _4339;
    assign _4342 = _1058 ? _4341 : _1001;
    assign _4338 = _1055 & _408;
    assign _4343 = _4338 ? _998 : _4342;
    assign _220 = _4343;
    always @(posedge _416) begin
        if (_414)
            _1001 <= _5492;
        else
            _1001 <= _220;
    end
    assign _1329 = { gnd,
                     _1001 };
    assign _1331 = _1329 < _1330;
    assign _4346 = _1331 ? _1001 : _998;
    assign _1323 = { gnd,
                     _995 };
    assign _1322 = { gnd,
                     _998 };
    assign _1324 = _1322 < _1323;
    assign _4345 = _1324 ? _995 : _998;
    assign _1321 = _1064[0:0];
    assign _4347 = _1321 ? _4346 : _4345;
    assign _4348 = _1058 ? _4347 : _998;
    assign _4344 = _1055 & _408;
    assign _4349 = _4344 ? _995 : _4348;
    assign _221 = _4349;
    always @(posedge _416) begin
        if (_414)
            _998 <= _5492;
        else
            _998 <= _221;
    end
    assign _1338 = { gnd,
                     _998 };
    assign _1340 = _1338 < _1339;
    assign _4351 = _1340 ? _998 : _995;
    assign _1337 = _1064[0:0];
    assign _4353 = _1337 ? _4352 : _4351;
    assign _4354 = _1058 ? _4353 : _995;
    assign _4350 = _1055 & _408;
    assign _4355 = _4350 ? _992 : _4354;
    assign _222 = _4355;
    always @(posedge _416) begin
        if (_414)
            _995 <= _5492;
        else
            _995 <= _222;
    end
    assign _1361 = { gnd,
                     _995 };
    assign _1363 = _1361 < _1362;
    assign _4358 = _1363 ? _995 : _992;
    assign _1355 = { gnd,
                     _989 };
    assign _1354 = { gnd,
                     _992 };
    assign _1356 = _1354 < _1355;
    assign _4357 = _1356 ? _989 : _992;
    assign _1353 = _1064[0:0];
    assign _4359 = _1353 ? _4358 : _4357;
    assign _4360 = _1058 ? _4359 : _992;
    assign _4356 = _1055 & _408;
    assign _4361 = _4356 ? _989 : _4360;
    assign _223 = _4361;
    always @(posedge _416) begin
        if (_414)
            _992 <= _5492;
        else
            _992 <= _223;
    end
    assign _1370 = { gnd,
                     _992 };
    assign _1372 = _1370 < _1371;
    assign _4363 = _1372 ? _992 : _989;
    assign _1369 = _1064[0:0];
    assign _4365 = _1369 ? _4364 : _4363;
    assign _4366 = _1058 ? _4365 : _989;
    assign _4362 = _1055 & _408;
    assign _4367 = _4362 ? _986 : _4366;
    assign _224 = _4367;
    always @(posedge _416) begin
        if (_414)
            _989 <= _5492;
        else
            _989 <= _224;
    end
    assign _1393 = { gnd,
                     _989 };
    assign _1395 = _1393 < _1394;
    assign _4370 = _1395 ? _989 : _986;
    assign _1387 = { gnd,
                     _983 };
    assign _1386 = { gnd,
                     _986 };
    assign _1388 = _1386 < _1387;
    assign _4369 = _1388 ? _983 : _986;
    assign _1385 = _1064[0:0];
    assign _4371 = _1385 ? _4370 : _4369;
    assign _4372 = _1058 ? _4371 : _986;
    assign _4368 = _1055 & _408;
    assign _4373 = _4368 ? _983 : _4372;
    assign _225 = _4373;
    always @(posedge _416) begin
        if (_414)
            _986 <= _5492;
        else
            _986 <= _225;
    end
    assign _1402 = { gnd,
                     _986 };
    assign _1404 = _1402 < _1403;
    assign _4375 = _1404 ? _986 : _983;
    assign _1401 = _1064[0:0];
    assign _4377 = _1401 ? _4376 : _4375;
    assign _4378 = _1058 ? _4377 : _983;
    assign _4374 = _1055 & _408;
    assign _4379 = _4374 ? _980 : _4378;
    assign _226 = _4379;
    always @(posedge _416) begin
        if (_414)
            _983 <= _5492;
        else
            _983 <= _226;
    end
    assign _1425 = { gnd,
                     _983 };
    assign _1427 = _1425 < _1426;
    assign _4382 = _1427 ? _983 : _980;
    assign _1419 = { gnd,
                     _977 };
    assign _1418 = { gnd,
                     _980 };
    assign _1420 = _1418 < _1419;
    assign _4381 = _1420 ? _977 : _980;
    assign _1417 = _1064[0:0];
    assign _4383 = _1417 ? _4382 : _4381;
    assign _4384 = _1058 ? _4383 : _980;
    assign _4380 = _1055 & _408;
    assign _4385 = _4380 ? _977 : _4384;
    assign _227 = _4385;
    always @(posedge _416) begin
        if (_414)
            _980 <= _5492;
        else
            _980 <= _227;
    end
    assign _1434 = { gnd,
                     _980 };
    assign _1436 = _1434 < _1435;
    assign _4387 = _1436 ? _980 : _977;
    assign _1433 = _1064[0:0];
    assign _4389 = _1433 ? _4388 : _4387;
    assign _4390 = _1058 ? _4389 : _977;
    assign _4386 = _1055 & _408;
    assign _4391 = _4386 ? _974 : _4390;
    assign _228 = _4391;
    always @(posedge _416) begin
        if (_414)
            _977 <= _5492;
        else
            _977 <= _228;
    end
    assign _1457 = { gnd,
                     _977 };
    assign _1459 = _1457 < _1458;
    assign _4394 = _1459 ? _977 : _974;
    assign _1451 = { gnd,
                     _971 };
    assign _1450 = { gnd,
                     _974 };
    assign _1452 = _1450 < _1451;
    assign _4393 = _1452 ? _971 : _974;
    assign _1449 = _1064[0:0];
    assign _4395 = _1449 ? _4394 : _4393;
    assign _4396 = _1058 ? _4395 : _974;
    assign _4392 = _1055 & _408;
    assign _4397 = _4392 ? _971 : _4396;
    assign _229 = _4397;
    always @(posedge _416) begin
        if (_414)
            _974 <= _5492;
        else
            _974 <= _229;
    end
    assign _1466 = { gnd,
                     _974 };
    assign _1468 = _1466 < _1467;
    assign _4399 = _1468 ? _974 : _971;
    assign _1465 = _1064[0:0];
    assign _4401 = _1465 ? _4400 : _4399;
    assign _4402 = _1058 ? _4401 : _971;
    assign _4398 = _1055 & _408;
    assign _4403 = _4398 ? _968 : _4402;
    assign _230 = _4403;
    always @(posedge _416) begin
        if (_414)
            _971 <= _5492;
        else
            _971 <= _230;
    end
    assign _1489 = { gnd,
                     _971 };
    assign _1491 = _1489 < _1490;
    assign _4406 = _1491 ? _971 : _968;
    assign _1483 = { gnd,
                     _965 };
    assign _1482 = { gnd,
                     _968 };
    assign _1484 = _1482 < _1483;
    assign _4405 = _1484 ? _965 : _968;
    assign _1481 = _1064[0:0];
    assign _4407 = _1481 ? _4406 : _4405;
    assign _4408 = _1058 ? _4407 : _968;
    assign _4404 = _1055 & _408;
    assign _4409 = _4404 ? _965 : _4408;
    assign _231 = _4409;
    always @(posedge _416) begin
        if (_414)
            _968 <= _5492;
        else
            _968 <= _231;
    end
    assign _1498 = { gnd,
                     _968 };
    assign _1500 = _1498 < _1499;
    assign _4411 = _1500 ? _968 : _965;
    assign _1497 = _1064[0:0];
    assign _4413 = _1497 ? _4412 : _4411;
    assign _4414 = _1058 ? _4413 : _965;
    assign _4410 = _1055 & _408;
    assign _4415 = _4410 ? _962 : _4414;
    assign _232 = _4415;
    always @(posedge _416) begin
        if (_414)
            _965 <= _5492;
        else
            _965 <= _232;
    end
    assign _1521 = { gnd,
                     _965 };
    assign _1523 = _1521 < _1522;
    assign _4418 = _1523 ? _965 : _962;
    assign _1515 = { gnd,
                     _959 };
    assign _1514 = { gnd,
                     _962 };
    assign _1516 = _1514 < _1515;
    assign _4417 = _1516 ? _959 : _962;
    assign _1513 = _1064[0:0];
    assign _4419 = _1513 ? _4418 : _4417;
    assign _4420 = _1058 ? _4419 : _962;
    assign _4416 = _1055 & _408;
    assign _4421 = _4416 ? _959 : _4420;
    assign _233 = _4421;
    always @(posedge _416) begin
        if (_414)
            _962 <= _5492;
        else
            _962 <= _233;
    end
    assign _1530 = { gnd,
                     _962 };
    assign _1532 = _1530 < _1531;
    assign _4423 = _1532 ? _962 : _959;
    assign _1529 = _1064[0:0];
    assign _4425 = _1529 ? _4424 : _4423;
    assign _4426 = _1058 ? _4425 : _959;
    assign _4422 = _1055 & _408;
    assign _4427 = _4422 ? _956 : _4426;
    assign _234 = _4427;
    always @(posedge _416) begin
        if (_414)
            _959 <= _5492;
        else
            _959 <= _234;
    end
    assign _1553 = { gnd,
                     _959 };
    assign _1555 = _1553 < _1554;
    assign _4430 = _1555 ? _959 : _956;
    assign _1547 = { gnd,
                     _953 };
    assign _1546 = { gnd,
                     _956 };
    assign _1548 = _1546 < _1547;
    assign _4429 = _1548 ? _953 : _956;
    assign _1545 = _1064[0:0];
    assign _4431 = _1545 ? _4430 : _4429;
    assign _4432 = _1058 ? _4431 : _956;
    assign _4428 = _1055 & _408;
    assign _4433 = _4428 ? _953 : _4432;
    assign _235 = _4433;
    always @(posedge _416) begin
        if (_414)
            _956 <= _5492;
        else
            _956 <= _235;
    end
    assign _1562 = { gnd,
                     _956 };
    assign _1564 = _1562 < _1563;
    assign _4435 = _1564 ? _956 : _953;
    assign _1561 = _1064[0:0];
    assign _4437 = _1561 ? _4436 : _4435;
    assign _4438 = _1058 ? _4437 : _953;
    assign _4434 = _1055 & _408;
    assign _4439 = _4434 ? _950 : _4438;
    assign _236 = _4439;
    always @(posedge _416) begin
        if (_414)
            _953 <= _5492;
        else
            _953 <= _236;
    end
    assign _1585 = { gnd,
                     _953 };
    assign _1587 = _1585 < _1586;
    assign _4442 = _1587 ? _953 : _950;
    assign _1579 = { gnd,
                     _947 };
    assign _1578 = { gnd,
                     _950 };
    assign _1580 = _1578 < _1579;
    assign _4441 = _1580 ? _947 : _950;
    assign _1577 = _1064[0:0];
    assign _4443 = _1577 ? _4442 : _4441;
    assign _4444 = _1058 ? _4443 : _950;
    assign _4440 = _1055 & _408;
    assign _4445 = _4440 ? _947 : _4444;
    assign _237 = _4445;
    always @(posedge _416) begin
        if (_414)
            _950 <= _5492;
        else
            _950 <= _237;
    end
    assign _1594 = { gnd,
                     _950 };
    assign _1596 = _1594 < _1595;
    assign _4447 = _1596 ? _950 : _947;
    assign _1593 = _1064[0:0];
    assign _4449 = _1593 ? _4448 : _4447;
    assign _4450 = _1058 ? _4449 : _947;
    assign _4446 = _1055 & _408;
    assign _4451 = _4446 ? _944 : _4450;
    assign _238 = _4451;
    always @(posedge _416) begin
        if (_414)
            _947 <= _5492;
        else
            _947 <= _238;
    end
    assign _1617 = { gnd,
                     _947 };
    assign _1619 = _1617 < _1618;
    assign _4454 = _1619 ? _947 : _944;
    assign _1611 = { gnd,
                     _941 };
    assign _1610 = { gnd,
                     _944 };
    assign _1612 = _1610 < _1611;
    assign _4453 = _1612 ? _941 : _944;
    assign _1609 = _1064[0:0];
    assign _4455 = _1609 ? _4454 : _4453;
    assign _4456 = _1058 ? _4455 : _944;
    assign _4452 = _1055 & _408;
    assign _4457 = _4452 ? _941 : _4456;
    assign _239 = _4457;
    always @(posedge _416) begin
        if (_414)
            _944 <= _5492;
        else
            _944 <= _239;
    end
    assign _1626 = { gnd,
                     _944 };
    assign _1628 = _1626 < _1627;
    assign _4459 = _1628 ? _944 : _941;
    assign _1625 = _1064[0:0];
    assign _4461 = _1625 ? _4460 : _4459;
    assign _4462 = _1058 ? _4461 : _941;
    assign _4458 = _1055 & _408;
    assign _4463 = _4458 ? _938 : _4462;
    assign _240 = _4463;
    always @(posedge _416) begin
        if (_414)
            _941 <= _5492;
        else
            _941 <= _240;
    end
    assign _1649 = { gnd,
                     _941 };
    assign _1651 = _1649 < _1650;
    assign _4466 = _1651 ? _941 : _938;
    assign _1643 = { gnd,
                     _935 };
    assign _1642 = { gnd,
                     _938 };
    assign _1644 = _1642 < _1643;
    assign _4465 = _1644 ? _935 : _938;
    assign _1641 = _1064[0:0];
    assign _4467 = _1641 ? _4466 : _4465;
    assign _4468 = _1058 ? _4467 : _938;
    assign _4464 = _1055 & _408;
    assign _4469 = _4464 ? _935 : _4468;
    assign _241 = _4469;
    always @(posedge _416) begin
        if (_414)
            _938 <= _5492;
        else
            _938 <= _241;
    end
    assign _1658 = { gnd,
                     _938 };
    assign _1660 = _1658 < _1659;
    assign _4471 = _1660 ? _938 : _935;
    assign _1657 = _1064[0:0];
    assign _4473 = _1657 ? _4472 : _4471;
    assign _4474 = _1058 ? _4473 : _935;
    assign _4470 = _1055 & _408;
    assign _4475 = _4470 ? _932 : _4474;
    assign _242 = _4475;
    always @(posedge _416) begin
        if (_414)
            _935 <= _5492;
        else
            _935 <= _242;
    end
    assign _1681 = { gnd,
                     _935 };
    assign _1683 = _1681 < _1682;
    assign _4478 = _1683 ? _935 : _932;
    assign _1675 = { gnd,
                     _929 };
    assign _1674 = { gnd,
                     _932 };
    assign _1676 = _1674 < _1675;
    assign _4477 = _1676 ? _929 : _932;
    assign _1673 = _1064[0:0];
    assign _4479 = _1673 ? _4478 : _4477;
    assign _4480 = _1058 ? _4479 : _932;
    assign _4476 = _1055 & _408;
    assign _4481 = _4476 ? _929 : _4480;
    assign _243 = _4481;
    always @(posedge _416) begin
        if (_414)
            _932 <= _5492;
        else
            _932 <= _243;
    end
    assign _1690 = { gnd,
                     _932 };
    assign _1692 = _1690 < _1691;
    assign _4483 = _1692 ? _932 : _929;
    assign _1689 = _1064[0:0];
    assign _4485 = _1689 ? _4484 : _4483;
    assign _4486 = _1058 ? _4485 : _929;
    assign _4482 = _1055 & _408;
    assign _4487 = _4482 ? _926 : _4486;
    assign _244 = _4487;
    always @(posedge _416) begin
        if (_414)
            _929 <= _5492;
        else
            _929 <= _244;
    end
    assign _1713 = { gnd,
                     _929 };
    assign _1715 = _1713 < _1714;
    assign _4490 = _1715 ? _929 : _926;
    assign _1707 = { gnd,
                     _923 };
    assign _1706 = { gnd,
                     _926 };
    assign _1708 = _1706 < _1707;
    assign _4489 = _1708 ? _923 : _926;
    assign _1705 = _1064[0:0];
    assign _4491 = _1705 ? _4490 : _4489;
    assign _4492 = _1058 ? _4491 : _926;
    assign _4488 = _1055 & _408;
    assign _4493 = _4488 ? _923 : _4492;
    assign _245 = _4493;
    always @(posedge _416) begin
        if (_414)
            _926 <= _5492;
        else
            _926 <= _245;
    end
    assign _1722 = { gnd,
                     _926 };
    assign _1724 = _1722 < _1723;
    assign _4495 = _1724 ? _926 : _923;
    assign _1721 = _1064[0:0];
    assign _4497 = _1721 ? _4496 : _4495;
    assign _4498 = _1058 ? _4497 : _923;
    assign _4494 = _1055 & _408;
    assign _4499 = _4494 ? _920 : _4498;
    assign _246 = _4499;
    always @(posedge _416) begin
        if (_414)
            _923 <= _5492;
        else
            _923 <= _246;
    end
    assign _1745 = { gnd,
                     _923 };
    assign _1747 = _1745 < _1746;
    assign _4502 = _1747 ? _923 : _920;
    assign _1739 = { gnd,
                     _917 };
    assign _1738 = { gnd,
                     _920 };
    assign _1740 = _1738 < _1739;
    assign _4501 = _1740 ? _917 : _920;
    assign _1737 = _1064[0:0];
    assign _4503 = _1737 ? _4502 : _4501;
    assign _4504 = _1058 ? _4503 : _920;
    assign _4500 = _1055 & _408;
    assign _4505 = _4500 ? _917 : _4504;
    assign _247 = _4505;
    always @(posedge _416) begin
        if (_414)
            _920 <= _5492;
        else
            _920 <= _247;
    end
    assign _1754 = { gnd,
                     _920 };
    assign _1756 = _1754 < _1755;
    assign _4507 = _1756 ? _920 : _917;
    assign _1753 = _1064[0:0];
    assign _4509 = _1753 ? _4508 : _4507;
    assign _4510 = _1058 ? _4509 : _917;
    assign _4506 = _1055 & _408;
    assign _4511 = _4506 ? _914 : _4510;
    assign _248 = _4511;
    always @(posedge _416) begin
        if (_414)
            _917 <= _5492;
        else
            _917 <= _248;
    end
    assign _1777 = { gnd,
                     _917 };
    assign _1779 = _1777 < _1778;
    assign _4514 = _1779 ? _917 : _914;
    assign _1771 = { gnd,
                     _911 };
    assign _1770 = { gnd,
                     _914 };
    assign _1772 = _1770 < _1771;
    assign _4513 = _1772 ? _911 : _914;
    assign _1769 = _1064[0:0];
    assign _4515 = _1769 ? _4514 : _4513;
    assign _4516 = _1058 ? _4515 : _914;
    assign _4512 = _1055 & _408;
    assign _4517 = _4512 ? _911 : _4516;
    assign _249 = _4517;
    always @(posedge _416) begin
        if (_414)
            _914 <= _5492;
        else
            _914 <= _249;
    end
    assign _1786 = { gnd,
                     _914 };
    assign _1788 = _1786 < _1787;
    assign _4519 = _1788 ? _914 : _911;
    assign _1785 = _1064[0:0];
    assign _4521 = _1785 ? _4520 : _4519;
    assign _4522 = _1058 ? _4521 : _911;
    assign _4518 = _1055 & _408;
    assign _4523 = _4518 ? _908 : _4522;
    assign _250 = _4523;
    always @(posedge _416) begin
        if (_414)
            _911 <= _5492;
        else
            _911 <= _250;
    end
    assign _1809 = { gnd,
                     _911 };
    assign _1811 = _1809 < _1810;
    assign _4526 = _1811 ? _911 : _908;
    assign _1803 = { gnd,
                     _905 };
    assign _1802 = { gnd,
                     _908 };
    assign _1804 = _1802 < _1803;
    assign _4525 = _1804 ? _905 : _908;
    assign _1801 = _1064[0:0];
    assign _4527 = _1801 ? _4526 : _4525;
    assign _4528 = _1058 ? _4527 : _908;
    assign _4524 = _1055 & _408;
    assign _4529 = _4524 ? _905 : _4528;
    assign _251 = _4529;
    always @(posedge _416) begin
        if (_414)
            _908 <= _5492;
        else
            _908 <= _251;
    end
    assign _1818 = { gnd,
                     _908 };
    assign _1820 = _1818 < _1819;
    assign _4531 = _1820 ? _908 : _905;
    assign _1817 = _1064[0:0];
    assign _4533 = _1817 ? _4532 : _4531;
    assign _4534 = _1058 ? _4533 : _905;
    assign _4530 = _1055 & _408;
    assign _4535 = _4530 ? _902 : _4534;
    assign _252 = _4535;
    always @(posedge _416) begin
        if (_414)
            _905 <= _5492;
        else
            _905 <= _252;
    end
    assign _1841 = { gnd,
                     _905 };
    assign _1843 = _1841 < _1842;
    assign _4538 = _1843 ? _905 : _902;
    assign _1835 = { gnd,
                     _899 };
    assign _1834 = { gnd,
                     _902 };
    assign _1836 = _1834 < _1835;
    assign _4537 = _1836 ? _899 : _902;
    assign _1833 = _1064[0:0];
    assign _4539 = _1833 ? _4538 : _4537;
    assign _4540 = _1058 ? _4539 : _902;
    assign _4536 = _1055 & _408;
    assign _4541 = _4536 ? _899 : _4540;
    assign _253 = _4541;
    always @(posedge _416) begin
        if (_414)
            _902 <= _5492;
        else
            _902 <= _253;
    end
    assign _1850 = { gnd,
                     _902 };
    assign _1852 = _1850 < _1851;
    assign _4543 = _1852 ? _902 : _899;
    assign _1849 = _1064[0:0];
    assign _4545 = _1849 ? _4544 : _4543;
    assign _4546 = _1058 ? _4545 : _899;
    assign _4542 = _1055 & _408;
    assign _4547 = _4542 ? _896 : _4546;
    assign _254 = _4547;
    always @(posedge _416) begin
        if (_414)
            _899 <= _5492;
        else
            _899 <= _254;
    end
    assign _1873 = { gnd,
                     _899 };
    assign _1875 = _1873 < _1874;
    assign _4550 = _1875 ? _899 : _896;
    assign _1867 = { gnd,
                     _893 };
    assign _1866 = { gnd,
                     _896 };
    assign _1868 = _1866 < _1867;
    assign _4549 = _1868 ? _893 : _896;
    assign _1865 = _1064[0:0];
    assign _4551 = _1865 ? _4550 : _4549;
    assign _4552 = _1058 ? _4551 : _896;
    assign _4548 = _1055 & _408;
    assign _4553 = _4548 ? _893 : _4552;
    assign _255 = _4553;
    always @(posedge _416) begin
        if (_414)
            _896 <= _5492;
        else
            _896 <= _255;
    end
    assign _1882 = { gnd,
                     _896 };
    assign _1884 = _1882 < _1883;
    assign _4555 = _1884 ? _896 : _893;
    assign _1881 = _1064[0:0];
    assign _4557 = _1881 ? _4556 : _4555;
    assign _4558 = _1058 ? _4557 : _893;
    assign _4554 = _1055 & _408;
    assign _4559 = _4554 ? _890 : _4558;
    assign _256 = _4559;
    always @(posedge _416) begin
        if (_414)
            _893 <= _5492;
        else
            _893 <= _256;
    end
    assign _1905 = { gnd,
                     _893 };
    assign _1907 = _1905 < _1906;
    assign _4562 = _1907 ? _893 : _890;
    assign _1899 = { gnd,
                     _887 };
    assign _1898 = { gnd,
                     _890 };
    assign _1900 = _1898 < _1899;
    assign _4561 = _1900 ? _887 : _890;
    assign _1897 = _1064[0:0];
    assign _4563 = _1897 ? _4562 : _4561;
    assign _4564 = _1058 ? _4563 : _890;
    assign _4560 = _1055 & _408;
    assign _4565 = _4560 ? _887 : _4564;
    assign _257 = _4565;
    always @(posedge _416) begin
        if (_414)
            _890 <= _5492;
        else
            _890 <= _257;
    end
    assign _1914 = { gnd,
                     _890 };
    assign _1916 = _1914 < _1915;
    assign _4567 = _1916 ? _890 : _887;
    assign _1913 = _1064[0:0];
    assign _4569 = _1913 ? _4568 : _4567;
    assign _4570 = _1058 ? _4569 : _887;
    assign _4566 = _1055 & _408;
    assign _4571 = _4566 ? _884 : _4570;
    assign _258 = _4571;
    always @(posedge _416) begin
        if (_414)
            _887 <= _5492;
        else
            _887 <= _258;
    end
    assign _1937 = { gnd,
                     _887 };
    assign _1939 = _1937 < _1938;
    assign _4574 = _1939 ? _887 : _884;
    assign _1931 = { gnd,
                     _881 };
    assign _1930 = { gnd,
                     _884 };
    assign _1932 = _1930 < _1931;
    assign _4573 = _1932 ? _881 : _884;
    assign _1929 = _1064[0:0];
    assign _4575 = _1929 ? _4574 : _4573;
    assign _4576 = _1058 ? _4575 : _884;
    assign _4572 = _1055 & _408;
    assign _4577 = _4572 ? _881 : _4576;
    assign _259 = _4577;
    always @(posedge _416) begin
        if (_414)
            _884 <= _5492;
        else
            _884 <= _259;
    end
    assign _1946 = { gnd,
                     _884 };
    assign _1948 = _1946 < _1947;
    assign _4579 = _1948 ? _884 : _881;
    assign _1945 = _1064[0:0];
    assign _4581 = _1945 ? _4580 : _4579;
    assign _4582 = _1058 ? _4581 : _881;
    assign _4578 = _1055 & _408;
    assign _4583 = _4578 ? _878 : _4582;
    assign _260 = _4583;
    always @(posedge _416) begin
        if (_414)
            _881 <= _5492;
        else
            _881 <= _260;
    end
    assign _1969 = { gnd,
                     _881 };
    assign _1971 = _1969 < _1970;
    assign _4586 = _1971 ? _881 : _878;
    assign _1963 = { gnd,
                     _875 };
    assign _1962 = { gnd,
                     _878 };
    assign _1964 = _1962 < _1963;
    assign _4585 = _1964 ? _875 : _878;
    assign _1961 = _1064[0:0];
    assign _4587 = _1961 ? _4586 : _4585;
    assign _4588 = _1058 ? _4587 : _878;
    assign _4584 = _1055 & _408;
    assign _4589 = _4584 ? _875 : _4588;
    assign _261 = _4589;
    always @(posedge _416) begin
        if (_414)
            _878 <= _5492;
        else
            _878 <= _261;
    end
    assign _1978 = { gnd,
                     _878 };
    assign _1980 = _1978 < _1979;
    assign _4591 = _1980 ? _878 : _875;
    assign _1977 = _1064[0:0];
    assign _4593 = _1977 ? _4592 : _4591;
    assign _4594 = _1058 ? _4593 : _875;
    assign _4590 = _1055 & _408;
    assign _4595 = _4590 ? _872 : _4594;
    assign _262 = _4595;
    always @(posedge _416) begin
        if (_414)
            _875 <= _5492;
        else
            _875 <= _262;
    end
    assign _2001 = { gnd,
                     _875 };
    assign _2003 = _2001 < _2002;
    assign _4598 = _2003 ? _875 : _872;
    assign _1995 = { gnd,
                     _869 };
    assign _1994 = { gnd,
                     _872 };
    assign _1996 = _1994 < _1995;
    assign _4597 = _1996 ? _869 : _872;
    assign _1993 = _1064[0:0];
    assign _4599 = _1993 ? _4598 : _4597;
    assign _4600 = _1058 ? _4599 : _872;
    assign _4596 = _1055 & _408;
    assign _4601 = _4596 ? _869 : _4600;
    assign _263 = _4601;
    always @(posedge _416) begin
        if (_414)
            _872 <= _5492;
        else
            _872 <= _263;
    end
    assign _2010 = { gnd,
                     _872 };
    assign _2012 = _2010 < _2011;
    assign _4603 = _2012 ? _872 : _869;
    assign _2009 = _1064[0:0];
    assign _4605 = _2009 ? _4604 : _4603;
    assign _4606 = _1058 ? _4605 : _869;
    assign _4602 = _1055 & _408;
    assign _4607 = _4602 ? _866 : _4606;
    assign _264 = _4607;
    always @(posedge _416) begin
        if (_414)
            _869 <= _5492;
        else
            _869 <= _264;
    end
    assign _2033 = { gnd,
                     _869 };
    assign _2035 = _2033 < _2034;
    assign _4610 = _2035 ? _869 : _866;
    assign _2027 = { gnd,
                     _863 };
    assign _2026 = { gnd,
                     _866 };
    assign _2028 = _2026 < _2027;
    assign _4609 = _2028 ? _863 : _866;
    assign _2025 = _1064[0:0];
    assign _4611 = _2025 ? _4610 : _4609;
    assign _4612 = _1058 ? _4611 : _866;
    assign _4608 = _1055 & _408;
    assign _4613 = _4608 ? _863 : _4612;
    assign _265 = _4613;
    always @(posedge _416) begin
        if (_414)
            _866 <= _5492;
        else
            _866 <= _265;
    end
    assign _2042 = { gnd,
                     _866 };
    assign _2044 = _2042 < _2043;
    assign _4615 = _2044 ? _866 : _863;
    assign _2041 = _1064[0:0];
    assign _4617 = _2041 ? _4616 : _4615;
    assign _4618 = _1058 ? _4617 : _863;
    assign _4614 = _1055 & _408;
    assign _4619 = _4614 ? _860 : _4618;
    assign _266 = _4619;
    always @(posedge _416) begin
        if (_414)
            _863 <= _5492;
        else
            _863 <= _266;
    end
    assign _2065 = { gnd,
                     _863 };
    assign _2067 = _2065 < _2066;
    assign _4622 = _2067 ? _863 : _860;
    assign _2059 = { gnd,
                     _857 };
    assign _2058 = { gnd,
                     _860 };
    assign _2060 = _2058 < _2059;
    assign _4621 = _2060 ? _857 : _860;
    assign _2057 = _1064[0:0];
    assign _4623 = _2057 ? _4622 : _4621;
    assign _4624 = _1058 ? _4623 : _860;
    assign _4620 = _1055 & _408;
    assign _4625 = _4620 ? _857 : _4624;
    assign _267 = _4625;
    always @(posedge _416) begin
        if (_414)
            _860 <= _5492;
        else
            _860 <= _267;
    end
    assign _2074 = { gnd,
                     _860 };
    assign _2076 = _2074 < _2075;
    assign _4627 = _2076 ? _860 : _857;
    assign _2073 = _1064[0:0];
    assign _4629 = _2073 ? _4628 : _4627;
    assign _4630 = _1058 ? _4629 : _857;
    assign _4626 = _1055 & _408;
    assign _4631 = _4626 ? _854 : _4630;
    assign _268 = _4631;
    always @(posedge _416) begin
        if (_414)
            _857 <= _5492;
        else
            _857 <= _268;
    end
    assign _2097 = { gnd,
                     _857 };
    assign _2099 = _2097 < _2098;
    assign _4634 = _2099 ? _857 : _854;
    assign _2091 = { gnd,
                     _851 };
    assign _2090 = { gnd,
                     _854 };
    assign _2092 = _2090 < _2091;
    assign _4633 = _2092 ? _851 : _854;
    assign _2089 = _1064[0:0];
    assign _4635 = _2089 ? _4634 : _4633;
    assign _4636 = _1058 ? _4635 : _854;
    assign _4632 = _1055 & _408;
    assign _4637 = _4632 ? _851 : _4636;
    assign _269 = _4637;
    always @(posedge _416) begin
        if (_414)
            _854 <= _5492;
        else
            _854 <= _269;
    end
    assign _2106 = { gnd,
                     _854 };
    assign _2108 = _2106 < _2107;
    assign _4639 = _2108 ? _854 : _851;
    assign _2105 = _1064[0:0];
    assign _4641 = _2105 ? _4640 : _4639;
    assign _4642 = _1058 ? _4641 : _851;
    assign _4638 = _1055 & _408;
    assign _4643 = _4638 ? _848 : _4642;
    assign _270 = _4643;
    always @(posedge _416) begin
        if (_414)
            _851 <= _5492;
        else
            _851 <= _270;
    end
    assign _2129 = { gnd,
                     _851 };
    assign _2131 = _2129 < _2130;
    assign _4646 = _2131 ? _851 : _848;
    assign _2123 = { gnd,
                     _845 };
    assign _2122 = { gnd,
                     _848 };
    assign _2124 = _2122 < _2123;
    assign _4645 = _2124 ? _845 : _848;
    assign _2121 = _1064[0:0];
    assign _4647 = _2121 ? _4646 : _4645;
    assign _4648 = _1058 ? _4647 : _848;
    assign _4644 = _1055 & _408;
    assign _4649 = _4644 ? _845 : _4648;
    assign _271 = _4649;
    always @(posedge _416) begin
        if (_414)
            _848 <= _5492;
        else
            _848 <= _271;
    end
    assign _2138 = { gnd,
                     _848 };
    assign _2140 = _2138 < _2139;
    assign _4651 = _2140 ? _848 : _845;
    assign _2137 = _1064[0:0];
    assign _4653 = _2137 ? _4652 : _4651;
    assign _4654 = _1058 ? _4653 : _845;
    assign _4650 = _1055 & _408;
    assign _4655 = _4650 ? _842 : _4654;
    assign _272 = _4655;
    always @(posedge _416) begin
        if (_414)
            _845 <= _5492;
        else
            _845 <= _272;
    end
    assign _2161 = { gnd,
                     _845 };
    assign _2163 = _2161 < _2162;
    assign _4658 = _2163 ? _845 : _842;
    assign _2155 = { gnd,
                     _839 };
    assign _2154 = { gnd,
                     _842 };
    assign _2156 = _2154 < _2155;
    assign _4657 = _2156 ? _839 : _842;
    assign _2153 = _1064[0:0];
    assign _4659 = _2153 ? _4658 : _4657;
    assign _4660 = _1058 ? _4659 : _842;
    assign _4656 = _1055 & _408;
    assign _4661 = _4656 ? _839 : _4660;
    assign _273 = _4661;
    always @(posedge _416) begin
        if (_414)
            _842 <= _5492;
        else
            _842 <= _273;
    end
    assign _2170 = { gnd,
                     _842 };
    assign _2172 = _2170 < _2171;
    assign _4663 = _2172 ? _842 : _839;
    assign _2169 = _1064[0:0];
    assign _4665 = _2169 ? _4664 : _4663;
    assign _4666 = _1058 ? _4665 : _839;
    assign _4662 = _1055 & _408;
    assign _4667 = _4662 ? _836 : _4666;
    assign _274 = _4667;
    always @(posedge _416) begin
        if (_414)
            _839 <= _5492;
        else
            _839 <= _274;
    end
    assign _2193 = { gnd,
                     _839 };
    assign _2195 = _2193 < _2194;
    assign _4670 = _2195 ? _839 : _836;
    assign _2187 = { gnd,
                     _833 };
    assign _2186 = { gnd,
                     _836 };
    assign _2188 = _2186 < _2187;
    assign _4669 = _2188 ? _833 : _836;
    assign _2185 = _1064[0:0];
    assign _4671 = _2185 ? _4670 : _4669;
    assign _4672 = _1058 ? _4671 : _836;
    assign _4668 = _1055 & _408;
    assign _4673 = _4668 ? _833 : _4672;
    assign _275 = _4673;
    always @(posedge _416) begin
        if (_414)
            _836 <= _5492;
        else
            _836 <= _275;
    end
    assign _2202 = { gnd,
                     _836 };
    assign _2204 = _2202 < _2203;
    assign _4675 = _2204 ? _836 : _833;
    assign _2201 = _1064[0:0];
    assign _4677 = _2201 ? _4676 : _4675;
    assign _4678 = _1058 ? _4677 : _833;
    assign _4674 = _1055 & _408;
    assign _4679 = _4674 ? _830 : _4678;
    assign _276 = _4679;
    always @(posedge _416) begin
        if (_414)
            _833 <= _5492;
        else
            _833 <= _276;
    end
    assign _2225 = { gnd,
                     _833 };
    assign _2227 = _2225 < _2226;
    assign _4682 = _2227 ? _833 : _830;
    assign _2219 = { gnd,
                     _827 };
    assign _2218 = { gnd,
                     _830 };
    assign _2220 = _2218 < _2219;
    assign _4681 = _2220 ? _827 : _830;
    assign _2217 = _1064[0:0];
    assign _4683 = _2217 ? _4682 : _4681;
    assign _4684 = _1058 ? _4683 : _830;
    assign _4680 = _1055 & _408;
    assign _4685 = _4680 ? _827 : _4684;
    assign _277 = _4685;
    always @(posedge _416) begin
        if (_414)
            _830 <= _5492;
        else
            _830 <= _277;
    end
    assign _2234 = { gnd,
                     _830 };
    assign _2236 = _2234 < _2235;
    assign _4687 = _2236 ? _830 : _827;
    assign _2233 = _1064[0:0];
    assign _4689 = _2233 ? _4688 : _4687;
    assign _4690 = _1058 ? _4689 : _827;
    assign _4686 = _1055 & _408;
    assign _4691 = _4686 ? _824 : _4690;
    assign _278 = _4691;
    always @(posedge _416) begin
        if (_414)
            _827 <= _5492;
        else
            _827 <= _278;
    end
    assign _2257 = { gnd,
                     _827 };
    assign _2259 = _2257 < _2258;
    assign _4694 = _2259 ? _827 : _824;
    assign _2251 = { gnd,
                     _821 };
    assign _2250 = { gnd,
                     _824 };
    assign _2252 = _2250 < _2251;
    assign _4693 = _2252 ? _821 : _824;
    assign _2249 = _1064[0:0];
    assign _4695 = _2249 ? _4694 : _4693;
    assign _4696 = _1058 ? _4695 : _824;
    assign _4692 = _1055 & _408;
    assign _4697 = _4692 ? _821 : _4696;
    assign _279 = _4697;
    always @(posedge _416) begin
        if (_414)
            _824 <= _5492;
        else
            _824 <= _279;
    end
    assign _2266 = { gnd,
                     _824 };
    assign _2268 = _2266 < _2267;
    assign _4699 = _2268 ? _824 : _821;
    assign _2265 = _1064[0:0];
    assign _4701 = _2265 ? _4700 : _4699;
    assign _4702 = _1058 ? _4701 : _821;
    assign _4698 = _1055 & _408;
    assign _4703 = _4698 ? _818 : _4702;
    assign _280 = _4703;
    always @(posedge _416) begin
        if (_414)
            _821 <= _5492;
        else
            _821 <= _280;
    end
    assign _2289 = { gnd,
                     _821 };
    assign _2291 = _2289 < _2290;
    assign _4706 = _2291 ? _821 : _818;
    assign _2283 = { gnd,
                     _815 };
    assign _2282 = { gnd,
                     _818 };
    assign _2284 = _2282 < _2283;
    assign _4705 = _2284 ? _815 : _818;
    assign _2281 = _1064[0:0];
    assign _4707 = _2281 ? _4706 : _4705;
    assign _4708 = _1058 ? _4707 : _818;
    assign _4704 = _1055 & _408;
    assign _4709 = _4704 ? _815 : _4708;
    assign _281 = _4709;
    always @(posedge _416) begin
        if (_414)
            _818 <= _5492;
        else
            _818 <= _281;
    end
    assign _2298 = { gnd,
                     _818 };
    assign _2300 = _2298 < _2299;
    assign _4711 = _2300 ? _818 : _815;
    assign _2297 = _1064[0:0];
    assign _4713 = _2297 ? _4712 : _4711;
    assign _4714 = _1058 ? _4713 : _815;
    assign _4710 = _1055 & _408;
    assign _4715 = _4710 ? _812 : _4714;
    assign _282 = _4715;
    always @(posedge _416) begin
        if (_414)
            _815 <= _5492;
        else
            _815 <= _282;
    end
    assign _2321 = { gnd,
                     _815 };
    assign _2323 = _2321 < _2322;
    assign _4718 = _2323 ? _815 : _812;
    assign _2315 = { gnd,
                     _809 };
    assign _2314 = { gnd,
                     _812 };
    assign _2316 = _2314 < _2315;
    assign _4717 = _2316 ? _809 : _812;
    assign _2313 = _1064[0:0];
    assign _4719 = _2313 ? _4718 : _4717;
    assign _4720 = _1058 ? _4719 : _812;
    assign _4716 = _1055 & _408;
    assign _4721 = _4716 ? _809 : _4720;
    assign _283 = _4721;
    always @(posedge _416) begin
        if (_414)
            _812 <= _5492;
        else
            _812 <= _283;
    end
    assign _2330 = { gnd,
                     _812 };
    assign _2332 = _2330 < _2331;
    assign _4723 = _2332 ? _812 : _809;
    assign _2329 = _1064[0:0];
    assign _4725 = _2329 ? _4724 : _4723;
    assign _4726 = _1058 ? _4725 : _809;
    assign _4722 = _1055 & _408;
    assign _4727 = _4722 ? _806 : _4726;
    assign _284 = _4727;
    always @(posedge _416) begin
        if (_414)
            _809 <= _5492;
        else
            _809 <= _284;
    end
    assign _2353 = { gnd,
                     _809 };
    assign _2355 = _2353 < _2354;
    assign _4730 = _2355 ? _809 : _806;
    assign _2347 = { gnd,
                     _803 };
    assign _2346 = { gnd,
                     _806 };
    assign _2348 = _2346 < _2347;
    assign _4729 = _2348 ? _803 : _806;
    assign _2345 = _1064[0:0];
    assign _4731 = _2345 ? _4730 : _4729;
    assign _4732 = _1058 ? _4731 : _806;
    assign _4728 = _1055 & _408;
    assign _4733 = _4728 ? _803 : _4732;
    assign _285 = _4733;
    always @(posedge _416) begin
        if (_414)
            _806 <= _5492;
        else
            _806 <= _285;
    end
    assign _2362 = { gnd,
                     _806 };
    assign _2364 = _2362 < _2363;
    assign _4735 = _2364 ? _806 : _803;
    assign _2361 = _1064[0:0];
    assign _4737 = _2361 ? _4736 : _4735;
    assign _4738 = _1058 ? _4737 : _803;
    assign _4734 = _1055 & _408;
    assign _4739 = _4734 ? _800 : _4738;
    assign _286 = _4739;
    always @(posedge _416) begin
        if (_414)
            _803 <= _5492;
        else
            _803 <= _286;
    end
    assign _2385 = { gnd,
                     _803 };
    assign _2387 = _2385 < _2386;
    assign _4742 = _2387 ? _803 : _800;
    assign _2379 = { gnd,
                     _797 };
    assign _2378 = { gnd,
                     _800 };
    assign _2380 = _2378 < _2379;
    assign _4741 = _2380 ? _797 : _800;
    assign _2377 = _1064[0:0];
    assign _4743 = _2377 ? _4742 : _4741;
    assign _4744 = _1058 ? _4743 : _800;
    assign _4740 = _1055 & _408;
    assign _4745 = _4740 ? _797 : _4744;
    assign _287 = _4745;
    always @(posedge _416) begin
        if (_414)
            _800 <= _5492;
        else
            _800 <= _287;
    end
    assign _2394 = { gnd,
                     _800 };
    assign _2396 = _2394 < _2395;
    assign _4747 = _2396 ? _800 : _797;
    assign _2393 = _1064[0:0];
    assign _4749 = _2393 ? _4748 : _4747;
    assign _4750 = _1058 ? _4749 : _797;
    assign _4746 = _1055 & _408;
    assign _4751 = _4746 ? _794 : _4750;
    assign _288 = _4751;
    always @(posedge _416) begin
        if (_414)
            _797 <= _5492;
        else
            _797 <= _288;
    end
    assign _2417 = { gnd,
                     _797 };
    assign _2419 = _2417 < _2418;
    assign _4754 = _2419 ? _797 : _794;
    assign _2411 = { gnd,
                     _791 };
    assign _2410 = { gnd,
                     _794 };
    assign _2412 = _2410 < _2411;
    assign _4753 = _2412 ? _791 : _794;
    assign _2409 = _1064[0:0];
    assign _4755 = _2409 ? _4754 : _4753;
    assign _4756 = _1058 ? _4755 : _794;
    assign _4752 = _1055 & _408;
    assign _4757 = _4752 ? _791 : _4756;
    assign _289 = _4757;
    always @(posedge _416) begin
        if (_414)
            _794 <= _5492;
        else
            _794 <= _289;
    end
    assign _2426 = { gnd,
                     _794 };
    assign _2428 = _2426 < _2427;
    assign _4759 = _2428 ? _794 : _791;
    assign _2425 = _1064[0:0];
    assign _4761 = _2425 ? _4760 : _4759;
    assign _4762 = _1058 ? _4761 : _791;
    assign _4758 = _1055 & _408;
    assign _4763 = _4758 ? _788 : _4762;
    assign _290 = _4763;
    always @(posedge _416) begin
        if (_414)
            _791 <= _5492;
        else
            _791 <= _290;
    end
    assign _2449 = { gnd,
                     _791 };
    assign _2451 = _2449 < _2450;
    assign _4766 = _2451 ? _791 : _788;
    assign _2443 = { gnd,
                     _785 };
    assign _2442 = { gnd,
                     _788 };
    assign _2444 = _2442 < _2443;
    assign _4765 = _2444 ? _785 : _788;
    assign _2441 = _1064[0:0];
    assign _4767 = _2441 ? _4766 : _4765;
    assign _4768 = _1058 ? _4767 : _788;
    assign _4764 = _1055 & _408;
    assign _4769 = _4764 ? _785 : _4768;
    assign _291 = _4769;
    always @(posedge _416) begin
        if (_414)
            _788 <= _5492;
        else
            _788 <= _291;
    end
    assign _2458 = { gnd,
                     _788 };
    assign _2460 = _2458 < _2459;
    assign _4771 = _2460 ? _788 : _785;
    assign _2457 = _1064[0:0];
    assign _4773 = _2457 ? _4772 : _4771;
    assign _4774 = _1058 ? _4773 : _785;
    assign _4770 = _1055 & _408;
    assign _4775 = _4770 ? _782 : _4774;
    assign _292 = _4775;
    always @(posedge _416) begin
        if (_414)
            _785 <= _5492;
        else
            _785 <= _292;
    end
    assign _2481 = { gnd,
                     _785 };
    assign _2483 = _2481 < _2482;
    assign _4778 = _2483 ? _785 : _782;
    assign _2475 = { gnd,
                     _779 };
    assign _2474 = { gnd,
                     _782 };
    assign _2476 = _2474 < _2475;
    assign _4777 = _2476 ? _779 : _782;
    assign _2473 = _1064[0:0];
    assign _4779 = _2473 ? _4778 : _4777;
    assign _4780 = _1058 ? _4779 : _782;
    assign _4776 = _1055 & _408;
    assign _4781 = _4776 ? _779 : _4780;
    assign _293 = _4781;
    always @(posedge _416) begin
        if (_414)
            _782 <= _5492;
        else
            _782 <= _293;
    end
    assign _2490 = { gnd,
                     _782 };
    assign _2492 = _2490 < _2491;
    assign _4783 = _2492 ? _782 : _779;
    assign _2489 = _1064[0:0];
    assign _4785 = _2489 ? _4784 : _4783;
    assign _4786 = _1058 ? _4785 : _779;
    assign _4782 = _1055 & _408;
    assign _4787 = _4782 ? _776 : _4786;
    assign _294 = _4787;
    always @(posedge _416) begin
        if (_414)
            _779 <= _5492;
        else
            _779 <= _294;
    end
    assign _2513 = { gnd,
                     _779 };
    assign _2515 = _2513 < _2514;
    assign _4790 = _2515 ? _779 : _776;
    assign _2507 = { gnd,
                     _773 };
    assign _2506 = { gnd,
                     _776 };
    assign _2508 = _2506 < _2507;
    assign _4789 = _2508 ? _773 : _776;
    assign _2505 = _1064[0:0];
    assign _4791 = _2505 ? _4790 : _4789;
    assign _4792 = _1058 ? _4791 : _776;
    assign _4788 = _1055 & _408;
    assign _4793 = _4788 ? _773 : _4792;
    assign _295 = _4793;
    always @(posedge _416) begin
        if (_414)
            _776 <= _5492;
        else
            _776 <= _295;
    end
    assign _2522 = { gnd,
                     _776 };
    assign _2524 = _2522 < _2523;
    assign _4795 = _2524 ? _776 : _773;
    assign _2521 = _1064[0:0];
    assign _4797 = _2521 ? _4796 : _4795;
    assign _4798 = _1058 ? _4797 : _773;
    assign _4794 = _1055 & _408;
    assign _4799 = _4794 ? _770 : _4798;
    assign _296 = _4799;
    always @(posedge _416) begin
        if (_414)
            _773 <= _5492;
        else
            _773 <= _296;
    end
    assign _2545 = { gnd,
                     _773 };
    assign _2547 = _2545 < _2546;
    assign _4802 = _2547 ? _773 : _770;
    assign _2539 = { gnd,
                     _767 };
    assign _2538 = { gnd,
                     _770 };
    assign _2540 = _2538 < _2539;
    assign _4801 = _2540 ? _767 : _770;
    assign _2537 = _1064[0:0];
    assign _4803 = _2537 ? _4802 : _4801;
    assign _4804 = _1058 ? _4803 : _770;
    assign _4800 = _1055 & _408;
    assign _4805 = _4800 ? _767 : _4804;
    assign _297 = _4805;
    always @(posedge _416) begin
        if (_414)
            _770 <= _5492;
        else
            _770 <= _297;
    end
    assign _2554 = { gnd,
                     _770 };
    assign _2556 = _2554 < _2555;
    assign _4807 = _2556 ? _770 : _767;
    assign _2553 = _1064[0:0];
    assign _4809 = _2553 ? _4808 : _4807;
    assign _4810 = _1058 ? _4809 : _767;
    assign _4806 = _1055 & _408;
    assign _4811 = _4806 ? _764 : _4810;
    assign _298 = _4811;
    always @(posedge _416) begin
        if (_414)
            _767 <= _5492;
        else
            _767 <= _298;
    end
    assign _2577 = { gnd,
                     _767 };
    assign _2579 = _2577 < _2578;
    assign _4814 = _2579 ? _767 : _764;
    assign _2571 = { gnd,
                     _761 };
    assign _2570 = { gnd,
                     _764 };
    assign _2572 = _2570 < _2571;
    assign _4813 = _2572 ? _761 : _764;
    assign _2569 = _1064[0:0];
    assign _4815 = _2569 ? _4814 : _4813;
    assign _4816 = _1058 ? _4815 : _764;
    assign _4812 = _1055 & _408;
    assign _4817 = _4812 ? _761 : _4816;
    assign _299 = _4817;
    always @(posedge _416) begin
        if (_414)
            _764 <= _5492;
        else
            _764 <= _299;
    end
    assign _2586 = { gnd,
                     _764 };
    assign _2588 = _2586 < _2587;
    assign _4819 = _2588 ? _764 : _761;
    assign _2585 = _1064[0:0];
    assign _4821 = _2585 ? _4820 : _4819;
    assign _4822 = _1058 ? _4821 : _761;
    assign _4818 = _1055 & _408;
    assign _4823 = _4818 ? _758 : _4822;
    assign _300 = _4823;
    always @(posedge _416) begin
        if (_414)
            _761 <= _5492;
        else
            _761 <= _300;
    end
    assign _2609 = { gnd,
                     _761 };
    assign _2611 = _2609 < _2610;
    assign _4826 = _2611 ? _761 : _758;
    assign _2603 = { gnd,
                     _755 };
    assign _2602 = { gnd,
                     _758 };
    assign _2604 = _2602 < _2603;
    assign _4825 = _2604 ? _755 : _758;
    assign _2601 = _1064[0:0];
    assign _4827 = _2601 ? _4826 : _4825;
    assign _4828 = _1058 ? _4827 : _758;
    assign _4824 = _1055 & _408;
    assign _4829 = _4824 ? _755 : _4828;
    assign _301 = _4829;
    always @(posedge _416) begin
        if (_414)
            _758 <= _5492;
        else
            _758 <= _301;
    end
    assign _2618 = { gnd,
                     _758 };
    assign _2620 = _2618 < _2619;
    assign _4831 = _2620 ? _758 : _755;
    assign _2617 = _1064[0:0];
    assign _4833 = _2617 ? _4832 : _4831;
    assign _4834 = _1058 ? _4833 : _755;
    assign _4830 = _1055 & _408;
    assign _4835 = _4830 ? _752 : _4834;
    assign _302 = _4835;
    always @(posedge _416) begin
        if (_414)
            _755 <= _5492;
        else
            _755 <= _302;
    end
    assign _2641 = { gnd,
                     _755 };
    assign _2643 = _2641 < _2642;
    assign _4838 = _2643 ? _755 : _752;
    assign _2635 = { gnd,
                     _749 };
    assign _2634 = { gnd,
                     _752 };
    assign _2636 = _2634 < _2635;
    assign _4837 = _2636 ? _749 : _752;
    assign _2633 = _1064[0:0];
    assign _4839 = _2633 ? _4838 : _4837;
    assign _4840 = _1058 ? _4839 : _752;
    assign _4836 = _1055 & _408;
    assign _4841 = _4836 ? _749 : _4840;
    assign _303 = _4841;
    always @(posedge _416) begin
        if (_414)
            _752 <= _5492;
        else
            _752 <= _303;
    end
    assign _2650 = { gnd,
                     _752 };
    assign _2652 = _2650 < _2651;
    assign _4843 = _2652 ? _752 : _749;
    assign _2649 = _1064[0:0];
    assign _4845 = _2649 ? _4844 : _4843;
    assign _4846 = _1058 ? _4845 : _749;
    assign _4842 = _1055 & _408;
    assign _4847 = _4842 ? _746 : _4846;
    assign _304 = _4847;
    always @(posedge _416) begin
        if (_414)
            _749 <= _5492;
        else
            _749 <= _304;
    end
    assign _2673 = { gnd,
                     _749 };
    assign _2675 = _2673 < _2674;
    assign _4850 = _2675 ? _749 : _746;
    assign _2667 = { gnd,
                     _743 };
    assign _2666 = { gnd,
                     _746 };
    assign _2668 = _2666 < _2667;
    assign _4849 = _2668 ? _743 : _746;
    assign _2665 = _1064[0:0];
    assign _4851 = _2665 ? _4850 : _4849;
    assign _4852 = _1058 ? _4851 : _746;
    assign _4848 = _1055 & _408;
    assign _4853 = _4848 ? _743 : _4852;
    assign _305 = _4853;
    always @(posedge _416) begin
        if (_414)
            _746 <= _5492;
        else
            _746 <= _305;
    end
    assign _2682 = { gnd,
                     _746 };
    assign _2684 = _2682 < _2683;
    assign _4855 = _2684 ? _746 : _743;
    assign _2681 = _1064[0:0];
    assign _4857 = _2681 ? _4856 : _4855;
    assign _4858 = _1058 ? _4857 : _743;
    assign _4854 = _1055 & _408;
    assign _4859 = _4854 ? _740 : _4858;
    assign _306 = _4859;
    always @(posedge _416) begin
        if (_414)
            _743 <= _5492;
        else
            _743 <= _306;
    end
    assign _2705 = { gnd,
                     _743 };
    assign _2707 = _2705 < _2706;
    assign _4862 = _2707 ? _743 : _740;
    assign _2699 = { gnd,
                     _737 };
    assign _2698 = { gnd,
                     _740 };
    assign _2700 = _2698 < _2699;
    assign _4861 = _2700 ? _737 : _740;
    assign _2697 = _1064[0:0];
    assign _4863 = _2697 ? _4862 : _4861;
    assign _4864 = _1058 ? _4863 : _740;
    assign _4860 = _1055 & _408;
    assign _4865 = _4860 ? _737 : _4864;
    assign _307 = _4865;
    always @(posedge _416) begin
        if (_414)
            _740 <= _5492;
        else
            _740 <= _307;
    end
    assign _2714 = { gnd,
                     _740 };
    assign _2716 = _2714 < _2715;
    assign _4867 = _2716 ? _740 : _737;
    assign _2713 = _1064[0:0];
    assign _4869 = _2713 ? _4868 : _4867;
    assign _4870 = _1058 ? _4869 : _737;
    assign _4866 = _1055 & _408;
    assign _4871 = _4866 ? _734 : _4870;
    assign _308 = _4871;
    always @(posedge _416) begin
        if (_414)
            _737 <= _5492;
        else
            _737 <= _308;
    end
    assign _2737 = { gnd,
                     _737 };
    assign _2739 = _2737 < _2738;
    assign _4874 = _2739 ? _737 : _734;
    assign _2731 = { gnd,
                     _731 };
    assign _2730 = { gnd,
                     _734 };
    assign _2732 = _2730 < _2731;
    assign _4873 = _2732 ? _731 : _734;
    assign _2729 = _1064[0:0];
    assign _4875 = _2729 ? _4874 : _4873;
    assign _4876 = _1058 ? _4875 : _734;
    assign _4872 = _1055 & _408;
    assign _4877 = _4872 ? _731 : _4876;
    assign _309 = _4877;
    always @(posedge _416) begin
        if (_414)
            _734 <= _5492;
        else
            _734 <= _309;
    end
    assign _2746 = { gnd,
                     _734 };
    assign _2748 = _2746 < _2747;
    assign _4879 = _2748 ? _734 : _731;
    assign _2745 = _1064[0:0];
    assign _4881 = _2745 ? _4880 : _4879;
    assign _4882 = _1058 ? _4881 : _731;
    assign _4878 = _1055 & _408;
    assign _4883 = _4878 ? _728 : _4882;
    assign _310 = _4883;
    always @(posedge _416) begin
        if (_414)
            _731 <= _5492;
        else
            _731 <= _310;
    end
    assign _2769 = { gnd,
                     _731 };
    assign _2771 = _2769 < _2770;
    assign _4886 = _2771 ? _731 : _728;
    assign _2763 = { gnd,
                     _725 };
    assign _2762 = { gnd,
                     _728 };
    assign _2764 = _2762 < _2763;
    assign _4885 = _2764 ? _725 : _728;
    assign _2761 = _1064[0:0];
    assign _4887 = _2761 ? _4886 : _4885;
    assign _4888 = _1058 ? _4887 : _728;
    assign _4884 = _1055 & _408;
    assign _4889 = _4884 ? _725 : _4888;
    assign _311 = _4889;
    always @(posedge _416) begin
        if (_414)
            _728 <= _5492;
        else
            _728 <= _311;
    end
    assign _2778 = { gnd,
                     _728 };
    assign _2780 = _2778 < _2779;
    assign _4891 = _2780 ? _728 : _725;
    assign _2777 = _1064[0:0];
    assign _4893 = _2777 ? _4892 : _4891;
    assign _4894 = _1058 ? _4893 : _725;
    assign _4890 = _1055 & _408;
    assign _4895 = _4890 ? _722 : _4894;
    assign _312 = _4895;
    always @(posedge _416) begin
        if (_414)
            _725 <= _5492;
        else
            _725 <= _312;
    end
    assign _2801 = { gnd,
                     _725 };
    assign _2803 = _2801 < _2802;
    assign _4898 = _2803 ? _725 : _722;
    assign _2795 = { gnd,
                     _719 };
    assign _2794 = { gnd,
                     _722 };
    assign _2796 = _2794 < _2795;
    assign _4897 = _2796 ? _719 : _722;
    assign _2793 = _1064[0:0];
    assign _4899 = _2793 ? _4898 : _4897;
    assign _4900 = _1058 ? _4899 : _722;
    assign _4896 = _1055 & _408;
    assign _4901 = _4896 ? _719 : _4900;
    assign _313 = _4901;
    always @(posedge _416) begin
        if (_414)
            _722 <= _5492;
        else
            _722 <= _313;
    end
    assign _2810 = { gnd,
                     _722 };
    assign _2812 = _2810 < _2811;
    assign _4903 = _2812 ? _722 : _719;
    assign _2809 = _1064[0:0];
    assign _4905 = _2809 ? _4904 : _4903;
    assign _4906 = _1058 ? _4905 : _719;
    assign _4902 = _1055 & _408;
    assign _4907 = _4902 ? _716 : _4906;
    assign _314 = _4907;
    always @(posedge _416) begin
        if (_414)
            _719 <= _5492;
        else
            _719 <= _314;
    end
    assign _2833 = { gnd,
                     _719 };
    assign _2835 = _2833 < _2834;
    assign _4910 = _2835 ? _719 : _716;
    assign _2827 = { gnd,
                     _713 };
    assign _2826 = { gnd,
                     _716 };
    assign _2828 = _2826 < _2827;
    assign _4909 = _2828 ? _713 : _716;
    assign _2825 = _1064[0:0];
    assign _4911 = _2825 ? _4910 : _4909;
    assign _4912 = _1058 ? _4911 : _716;
    assign _4908 = _1055 & _408;
    assign _4913 = _4908 ? _713 : _4912;
    assign _315 = _4913;
    always @(posedge _416) begin
        if (_414)
            _716 <= _5492;
        else
            _716 <= _315;
    end
    assign _2842 = { gnd,
                     _716 };
    assign _2844 = _2842 < _2843;
    assign _4915 = _2844 ? _716 : _713;
    assign _2841 = _1064[0:0];
    assign _4917 = _2841 ? _4916 : _4915;
    assign _4918 = _1058 ? _4917 : _713;
    assign _4914 = _1055 & _408;
    assign _4919 = _4914 ? _710 : _4918;
    assign _316 = _4919;
    always @(posedge _416) begin
        if (_414)
            _713 <= _5492;
        else
            _713 <= _316;
    end
    assign _2865 = { gnd,
                     _713 };
    assign _2867 = _2865 < _2866;
    assign _4922 = _2867 ? _713 : _710;
    assign _2859 = { gnd,
                     _707 };
    assign _2858 = { gnd,
                     _710 };
    assign _2860 = _2858 < _2859;
    assign _4921 = _2860 ? _707 : _710;
    assign _2857 = _1064[0:0];
    assign _4923 = _2857 ? _4922 : _4921;
    assign _4924 = _1058 ? _4923 : _710;
    assign _4920 = _1055 & _408;
    assign _4925 = _4920 ? _707 : _4924;
    assign _317 = _4925;
    always @(posedge _416) begin
        if (_414)
            _710 <= _5492;
        else
            _710 <= _317;
    end
    assign _2874 = { gnd,
                     _710 };
    assign _2876 = _2874 < _2875;
    assign _4927 = _2876 ? _710 : _707;
    assign _2873 = _1064[0:0];
    assign _4929 = _2873 ? _4928 : _4927;
    assign _4930 = _1058 ? _4929 : _707;
    assign _4926 = _1055 & _408;
    assign _4931 = _4926 ? _704 : _4930;
    assign _318 = _4931;
    always @(posedge _416) begin
        if (_414)
            _707 <= _5492;
        else
            _707 <= _318;
    end
    assign _2897 = { gnd,
                     _707 };
    assign _2899 = _2897 < _2898;
    assign _4934 = _2899 ? _707 : _704;
    assign _2891 = { gnd,
                     _701 };
    assign _2890 = { gnd,
                     _704 };
    assign _2892 = _2890 < _2891;
    assign _4933 = _2892 ? _701 : _704;
    assign _2889 = _1064[0:0];
    assign _4935 = _2889 ? _4934 : _4933;
    assign _4936 = _1058 ? _4935 : _704;
    assign _4932 = _1055 & _408;
    assign _4937 = _4932 ? _701 : _4936;
    assign _319 = _4937;
    always @(posedge _416) begin
        if (_414)
            _704 <= _5492;
        else
            _704 <= _319;
    end
    assign _2906 = { gnd,
                     _704 };
    assign _2908 = _2906 < _2907;
    assign _4939 = _2908 ? _704 : _701;
    assign _2905 = _1064[0:0];
    assign _4941 = _2905 ? _4940 : _4939;
    assign _4942 = _1058 ? _4941 : _701;
    assign _4938 = _1055 & _408;
    assign _4943 = _4938 ? _698 : _4942;
    assign _320 = _4943;
    always @(posedge _416) begin
        if (_414)
            _701 <= _5492;
        else
            _701 <= _320;
    end
    assign _2929 = { gnd,
                     _701 };
    assign _2931 = _2929 < _2930;
    assign _4946 = _2931 ? _701 : _698;
    assign _2923 = { gnd,
                     _695 };
    assign _2922 = { gnd,
                     _698 };
    assign _2924 = _2922 < _2923;
    assign _4945 = _2924 ? _695 : _698;
    assign _2921 = _1064[0:0];
    assign _4947 = _2921 ? _4946 : _4945;
    assign _4948 = _1058 ? _4947 : _698;
    assign _4944 = _1055 & _408;
    assign _4949 = _4944 ? _695 : _4948;
    assign _321 = _4949;
    always @(posedge _416) begin
        if (_414)
            _698 <= _5492;
        else
            _698 <= _321;
    end
    assign _2938 = { gnd,
                     _698 };
    assign _2940 = _2938 < _2939;
    assign _4951 = _2940 ? _698 : _695;
    assign _2937 = _1064[0:0];
    assign _4953 = _2937 ? _4952 : _4951;
    assign _4954 = _1058 ? _4953 : _695;
    assign _4950 = _1055 & _408;
    assign _4955 = _4950 ? _692 : _4954;
    assign _322 = _4955;
    always @(posedge _416) begin
        if (_414)
            _695 <= _5492;
        else
            _695 <= _322;
    end
    assign _2961 = { gnd,
                     _695 };
    assign _2963 = _2961 < _2962;
    assign _4958 = _2963 ? _695 : _692;
    assign _2955 = { gnd,
                     _689 };
    assign _2954 = { gnd,
                     _692 };
    assign _2956 = _2954 < _2955;
    assign _4957 = _2956 ? _689 : _692;
    assign _2953 = _1064[0:0];
    assign _4959 = _2953 ? _4958 : _4957;
    assign _4960 = _1058 ? _4959 : _692;
    assign _4956 = _1055 & _408;
    assign _4961 = _4956 ? _689 : _4960;
    assign _323 = _4961;
    always @(posedge _416) begin
        if (_414)
            _692 <= _5492;
        else
            _692 <= _323;
    end
    assign _2970 = { gnd,
                     _692 };
    assign _2972 = _2970 < _2971;
    assign _4963 = _2972 ? _692 : _689;
    assign _2969 = _1064[0:0];
    assign _4965 = _2969 ? _4964 : _4963;
    assign _4966 = _1058 ? _4965 : _689;
    assign _4962 = _1055 & _408;
    assign _4967 = _4962 ? _686 : _4966;
    assign _324 = _4967;
    always @(posedge _416) begin
        if (_414)
            _689 <= _5492;
        else
            _689 <= _324;
    end
    assign _2993 = { gnd,
                     _689 };
    assign _2995 = _2993 < _2994;
    assign _4970 = _2995 ? _689 : _686;
    assign _2987 = { gnd,
                     _683 };
    assign _2986 = { gnd,
                     _686 };
    assign _2988 = _2986 < _2987;
    assign _4969 = _2988 ? _683 : _686;
    assign _2985 = _1064[0:0];
    assign _4971 = _2985 ? _4970 : _4969;
    assign _4972 = _1058 ? _4971 : _686;
    assign _4968 = _1055 & _408;
    assign _4973 = _4968 ? _683 : _4972;
    assign _325 = _4973;
    always @(posedge _416) begin
        if (_414)
            _686 <= _5492;
        else
            _686 <= _325;
    end
    assign _3002 = { gnd,
                     _686 };
    assign _3004 = _3002 < _3003;
    assign _4975 = _3004 ? _686 : _683;
    assign _3001 = _1064[0:0];
    assign _4977 = _3001 ? _4976 : _4975;
    assign _4978 = _1058 ? _4977 : _683;
    assign _4974 = _1055 & _408;
    assign _4979 = _4974 ? _680 : _4978;
    assign _326 = _4979;
    always @(posedge _416) begin
        if (_414)
            _683 <= _5492;
        else
            _683 <= _326;
    end
    assign _3025 = { gnd,
                     _683 };
    assign _3027 = _3025 < _3026;
    assign _4982 = _3027 ? _683 : _680;
    assign _3019 = { gnd,
                     _677 };
    assign _3018 = { gnd,
                     _680 };
    assign _3020 = _3018 < _3019;
    assign _4981 = _3020 ? _677 : _680;
    assign _3017 = _1064[0:0];
    assign _4983 = _3017 ? _4982 : _4981;
    assign _4984 = _1058 ? _4983 : _680;
    assign _4980 = _1055 & _408;
    assign _4985 = _4980 ? _677 : _4984;
    assign _327 = _4985;
    always @(posedge _416) begin
        if (_414)
            _680 <= _5492;
        else
            _680 <= _327;
    end
    assign _3034 = { gnd,
                     _680 };
    assign _3036 = _3034 < _3035;
    assign _4987 = _3036 ? _680 : _677;
    assign _3033 = _1064[0:0];
    assign _4989 = _3033 ? _4988 : _4987;
    assign _4990 = _1058 ? _4989 : _677;
    assign _4986 = _1055 & _408;
    assign _4991 = _4986 ? _674 : _4990;
    assign _328 = _4991;
    always @(posedge _416) begin
        if (_414)
            _677 <= _5492;
        else
            _677 <= _328;
    end
    assign _3057 = { gnd,
                     _677 };
    assign _3059 = _3057 < _3058;
    assign _4994 = _3059 ? _677 : _674;
    assign _3051 = { gnd,
                     _671 };
    assign _3050 = { gnd,
                     _674 };
    assign _3052 = _3050 < _3051;
    assign _4993 = _3052 ? _671 : _674;
    assign _3049 = _1064[0:0];
    assign _4995 = _3049 ? _4994 : _4993;
    assign _4996 = _1058 ? _4995 : _674;
    assign _4992 = _1055 & _408;
    assign _4997 = _4992 ? _671 : _4996;
    assign _329 = _4997;
    always @(posedge _416) begin
        if (_414)
            _674 <= _5492;
        else
            _674 <= _329;
    end
    assign _3066 = { gnd,
                     _674 };
    assign _3068 = _3066 < _3067;
    assign _4999 = _3068 ? _674 : _671;
    assign _3065 = _1064[0:0];
    assign _5001 = _3065 ? _5000 : _4999;
    assign _5002 = _1058 ? _5001 : _671;
    assign _4998 = _1055 & _408;
    assign _5003 = _4998 ? _668 : _5002;
    assign _330 = _5003;
    always @(posedge _416) begin
        if (_414)
            _671 <= _5492;
        else
            _671 <= _330;
    end
    assign _3089 = { gnd,
                     _671 };
    assign _3091 = _3089 < _3090;
    assign _5006 = _3091 ? _671 : _668;
    assign _3083 = { gnd,
                     _665 };
    assign _3082 = { gnd,
                     _668 };
    assign _3084 = _3082 < _3083;
    assign _5005 = _3084 ? _665 : _668;
    assign _3081 = _1064[0:0];
    assign _5007 = _3081 ? _5006 : _5005;
    assign _5008 = _1058 ? _5007 : _668;
    assign _5004 = _1055 & _408;
    assign _5009 = _5004 ? _665 : _5008;
    assign _331 = _5009;
    always @(posedge _416) begin
        if (_414)
            _668 <= _5492;
        else
            _668 <= _331;
    end
    assign _3098 = { gnd,
                     _668 };
    assign _3100 = _3098 < _3099;
    assign _5011 = _3100 ? _668 : _665;
    assign _3097 = _1064[0:0];
    assign _5013 = _3097 ? _5012 : _5011;
    assign _5014 = _1058 ? _5013 : _665;
    assign _5010 = _1055 & _408;
    assign _5015 = _5010 ? _662 : _5014;
    assign _332 = _5015;
    always @(posedge _416) begin
        if (_414)
            _665 <= _5492;
        else
            _665 <= _332;
    end
    assign _3121 = { gnd,
                     _665 };
    assign _3123 = _3121 < _3122;
    assign _5018 = _3123 ? _665 : _662;
    assign _3115 = { gnd,
                     _659 };
    assign _3114 = { gnd,
                     _662 };
    assign _3116 = _3114 < _3115;
    assign _5017 = _3116 ? _659 : _662;
    assign _3113 = _1064[0:0];
    assign _5019 = _3113 ? _5018 : _5017;
    assign _5020 = _1058 ? _5019 : _662;
    assign _5016 = _1055 & _408;
    assign _5021 = _5016 ? _659 : _5020;
    assign _333 = _5021;
    always @(posedge _416) begin
        if (_414)
            _662 <= _5492;
        else
            _662 <= _333;
    end
    assign _3130 = { gnd,
                     _662 };
    assign _3132 = _3130 < _3131;
    assign _5023 = _3132 ? _662 : _659;
    assign _3129 = _1064[0:0];
    assign _5025 = _3129 ? _5024 : _5023;
    assign _5026 = _1058 ? _5025 : _659;
    assign _5022 = _1055 & _408;
    assign _5027 = _5022 ? _656 : _5026;
    assign _334 = _5027;
    always @(posedge _416) begin
        if (_414)
            _659 <= _5492;
        else
            _659 <= _334;
    end
    assign _3153 = { gnd,
                     _659 };
    assign _3155 = _3153 < _3154;
    assign _5030 = _3155 ? _659 : _656;
    assign _3147 = { gnd,
                     _653 };
    assign _3146 = { gnd,
                     _656 };
    assign _3148 = _3146 < _3147;
    assign _5029 = _3148 ? _653 : _656;
    assign _3145 = _1064[0:0];
    assign _5031 = _3145 ? _5030 : _5029;
    assign _5032 = _1058 ? _5031 : _656;
    assign _5028 = _1055 & _408;
    assign _5033 = _5028 ? _653 : _5032;
    assign _335 = _5033;
    always @(posedge _416) begin
        if (_414)
            _656 <= _5492;
        else
            _656 <= _335;
    end
    assign _3162 = { gnd,
                     _656 };
    assign _3164 = _3162 < _3163;
    assign _5035 = _3164 ? _656 : _653;
    assign _3161 = _1064[0:0];
    assign _5037 = _3161 ? _5036 : _5035;
    assign _5038 = _1058 ? _5037 : _653;
    assign _5034 = _1055 & _408;
    assign _5039 = _5034 ? _650 : _5038;
    assign _336 = _5039;
    always @(posedge _416) begin
        if (_414)
            _653 <= _5492;
        else
            _653 <= _336;
    end
    assign _3185 = { gnd,
                     _653 };
    assign _3187 = _3185 < _3186;
    assign _5042 = _3187 ? _653 : _650;
    assign _3179 = { gnd,
                     _647 };
    assign _3178 = { gnd,
                     _650 };
    assign _3180 = _3178 < _3179;
    assign _5041 = _3180 ? _647 : _650;
    assign _3177 = _1064[0:0];
    assign _5043 = _3177 ? _5042 : _5041;
    assign _5044 = _1058 ? _5043 : _650;
    assign _5040 = _1055 & _408;
    assign _5045 = _5040 ? _647 : _5044;
    assign _337 = _5045;
    always @(posedge _416) begin
        if (_414)
            _650 <= _5492;
        else
            _650 <= _337;
    end
    assign _3194 = { gnd,
                     _650 };
    assign _3196 = _3194 < _3195;
    assign _5047 = _3196 ? _650 : _647;
    assign _3193 = _1064[0:0];
    assign _5049 = _3193 ? _5048 : _5047;
    assign _5050 = _1058 ? _5049 : _647;
    assign _5046 = _1055 & _408;
    assign _5051 = _5046 ? _644 : _5050;
    assign _338 = _5051;
    always @(posedge _416) begin
        if (_414)
            _647 <= _5492;
        else
            _647 <= _338;
    end
    assign _3217 = { gnd,
                     _647 };
    assign _3219 = _3217 < _3218;
    assign _5054 = _3219 ? _647 : _644;
    assign _3211 = { gnd,
                     _641 };
    assign _3210 = { gnd,
                     _644 };
    assign _3212 = _3210 < _3211;
    assign _5053 = _3212 ? _641 : _644;
    assign _3209 = _1064[0:0];
    assign _5055 = _3209 ? _5054 : _5053;
    assign _5056 = _1058 ? _5055 : _644;
    assign _5052 = _1055 & _408;
    assign _5057 = _5052 ? _641 : _5056;
    assign _339 = _5057;
    always @(posedge _416) begin
        if (_414)
            _644 <= _5492;
        else
            _644 <= _339;
    end
    assign _3226 = { gnd,
                     _644 };
    assign _3228 = _3226 < _3227;
    assign _5059 = _3228 ? _644 : _641;
    assign _3225 = _1064[0:0];
    assign _5061 = _3225 ? _5060 : _5059;
    assign _5062 = _1058 ? _5061 : _641;
    assign _5058 = _1055 & _408;
    assign _5063 = _5058 ? _638 : _5062;
    assign _340 = _5063;
    always @(posedge _416) begin
        if (_414)
            _641 <= _5492;
        else
            _641 <= _340;
    end
    assign _3249 = { gnd,
                     _641 };
    assign _3251 = _3249 < _3250;
    assign _5066 = _3251 ? _641 : _638;
    assign _3243 = { gnd,
                     _635 };
    assign _3242 = { gnd,
                     _638 };
    assign _3244 = _3242 < _3243;
    assign _5065 = _3244 ? _635 : _638;
    assign _3241 = _1064[0:0];
    assign _5067 = _3241 ? _5066 : _5065;
    assign _5068 = _1058 ? _5067 : _638;
    assign _5064 = _1055 & _408;
    assign _5069 = _5064 ? _635 : _5068;
    assign _341 = _5069;
    always @(posedge _416) begin
        if (_414)
            _638 <= _5492;
        else
            _638 <= _341;
    end
    assign _3258 = { gnd,
                     _638 };
    assign _3260 = _3258 < _3259;
    assign _5071 = _3260 ? _638 : _635;
    assign _3257 = _1064[0:0];
    assign _5073 = _3257 ? _5072 : _5071;
    assign _5074 = _1058 ? _5073 : _635;
    assign _5070 = _1055 & _408;
    assign _5075 = _5070 ? _632 : _5074;
    assign _342 = _5075;
    always @(posedge _416) begin
        if (_414)
            _635 <= _5492;
        else
            _635 <= _342;
    end
    assign _3281 = { gnd,
                     _635 };
    assign _3283 = _3281 < _3282;
    assign _5078 = _3283 ? _635 : _632;
    assign _3275 = { gnd,
                     _629 };
    assign _3274 = { gnd,
                     _632 };
    assign _3276 = _3274 < _3275;
    assign _5077 = _3276 ? _629 : _632;
    assign _3273 = _1064[0:0];
    assign _5079 = _3273 ? _5078 : _5077;
    assign _5080 = _1058 ? _5079 : _632;
    assign _5076 = _1055 & _408;
    assign _5081 = _5076 ? _629 : _5080;
    assign _343 = _5081;
    always @(posedge _416) begin
        if (_414)
            _632 <= _5492;
        else
            _632 <= _343;
    end
    assign _3290 = { gnd,
                     _632 };
    assign _3292 = _3290 < _3291;
    assign _5083 = _3292 ? _632 : _629;
    assign _3289 = _1064[0:0];
    assign _5085 = _3289 ? _5084 : _5083;
    assign _5086 = _1058 ? _5085 : _629;
    assign _5082 = _1055 & _408;
    assign _5087 = _5082 ? _626 : _5086;
    assign _344 = _5087;
    always @(posedge _416) begin
        if (_414)
            _629 <= _5492;
        else
            _629 <= _344;
    end
    assign _3313 = { gnd,
                     _629 };
    assign _3315 = _3313 < _3314;
    assign _5090 = _3315 ? _629 : _626;
    assign _3307 = { gnd,
                     _623 };
    assign _3306 = { gnd,
                     _626 };
    assign _3308 = _3306 < _3307;
    assign _5089 = _3308 ? _623 : _626;
    assign _3305 = _1064[0:0];
    assign _5091 = _3305 ? _5090 : _5089;
    assign _5092 = _1058 ? _5091 : _626;
    assign _5088 = _1055 & _408;
    assign _5093 = _5088 ? _623 : _5092;
    assign _345 = _5093;
    always @(posedge _416) begin
        if (_414)
            _626 <= _5492;
        else
            _626 <= _345;
    end
    assign _3322 = { gnd,
                     _626 };
    assign _3324 = _3322 < _3323;
    assign _5095 = _3324 ? _626 : _623;
    assign _3321 = _1064[0:0];
    assign _5097 = _3321 ? _5096 : _5095;
    assign _5098 = _1058 ? _5097 : _623;
    assign _5094 = _1055 & _408;
    assign _5099 = _5094 ? _620 : _5098;
    assign _346 = _5099;
    always @(posedge _416) begin
        if (_414)
            _623 <= _5492;
        else
            _623 <= _346;
    end
    assign _3345 = { gnd,
                     _623 };
    assign _3347 = _3345 < _3346;
    assign _5102 = _3347 ? _623 : _620;
    assign _3339 = { gnd,
                     _617 };
    assign _3338 = { gnd,
                     _620 };
    assign _3340 = _3338 < _3339;
    assign _5101 = _3340 ? _617 : _620;
    assign _3337 = _1064[0:0];
    assign _5103 = _3337 ? _5102 : _5101;
    assign _5104 = _1058 ? _5103 : _620;
    assign _5100 = _1055 & _408;
    assign _5105 = _5100 ? _617 : _5104;
    assign _347 = _5105;
    always @(posedge _416) begin
        if (_414)
            _620 <= _5492;
        else
            _620 <= _347;
    end
    assign _3354 = { gnd,
                     _620 };
    assign _3356 = _3354 < _3355;
    assign _5107 = _3356 ? _620 : _617;
    assign _3353 = _1064[0:0];
    assign _5109 = _3353 ? _5108 : _5107;
    assign _5110 = _1058 ? _5109 : _617;
    assign _5106 = _1055 & _408;
    assign _5111 = _5106 ? _614 : _5110;
    assign _348 = _5111;
    always @(posedge _416) begin
        if (_414)
            _617 <= _5492;
        else
            _617 <= _348;
    end
    assign _3377 = { gnd,
                     _617 };
    assign _3379 = _3377 < _3378;
    assign _5114 = _3379 ? _617 : _614;
    assign _3371 = { gnd,
                     _611 };
    assign _3370 = { gnd,
                     _614 };
    assign _3372 = _3370 < _3371;
    assign _5113 = _3372 ? _611 : _614;
    assign _3369 = _1064[0:0];
    assign _5115 = _3369 ? _5114 : _5113;
    assign _5116 = _1058 ? _5115 : _614;
    assign _5112 = _1055 & _408;
    assign _5117 = _5112 ? _611 : _5116;
    assign _349 = _5117;
    always @(posedge _416) begin
        if (_414)
            _614 <= _5492;
        else
            _614 <= _349;
    end
    assign _3386 = { gnd,
                     _614 };
    assign _3388 = _3386 < _3387;
    assign _5119 = _3388 ? _614 : _611;
    assign _3385 = _1064[0:0];
    assign _5121 = _3385 ? _5120 : _5119;
    assign _5122 = _1058 ? _5121 : _611;
    assign _5118 = _1055 & _408;
    assign _5123 = _5118 ? _608 : _5122;
    assign _350 = _5123;
    always @(posedge _416) begin
        if (_414)
            _611 <= _5492;
        else
            _611 <= _350;
    end
    assign _3409 = { gnd,
                     _611 };
    assign _3411 = _3409 < _3410;
    assign _5126 = _3411 ? _611 : _608;
    assign _3403 = { gnd,
                     _605 };
    assign _3402 = { gnd,
                     _608 };
    assign _3404 = _3402 < _3403;
    assign _5125 = _3404 ? _605 : _608;
    assign _3401 = _1064[0:0];
    assign _5127 = _3401 ? _5126 : _5125;
    assign _5128 = _1058 ? _5127 : _608;
    assign _5124 = _1055 & _408;
    assign _5129 = _5124 ? _605 : _5128;
    assign _351 = _5129;
    always @(posedge _416) begin
        if (_414)
            _608 <= _5492;
        else
            _608 <= _351;
    end
    assign _3418 = { gnd,
                     _608 };
    assign _3420 = _3418 < _3419;
    assign _5131 = _3420 ? _608 : _605;
    assign _3417 = _1064[0:0];
    assign _5133 = _3417 ? _5132 : _5131;
    assign _5134 = _1058 ? _5133 : _605;
    assign _5130 = _1055 & _408;
    assign _5135 = _5130 ? _602 : _5134;
    assign _352 = _5135;
    always @(posedge _416) begin
        if (_414)
            _605 <= _5492;
        else
            _605 <= _352;
    end
    assign _3441 = { gnd,
                     _605 };
    assign _3443 = _3441 < _3442;
    assign _5138 = _3443 ? _605 : _602;
    assign _3435 = { gnd,
                     _599 };
    assign _3434 = { gnd,
                     _602 };
    assign _3436 = _3434 < _3435;
    assign _5137 = _3436 ? _599 : _602;
    assign _3433 = _1064[0:0];
    assign _5139 = _3433 ? _5138 : _5137;
    assign _5140 = _1058 ? _5139 : _602;
    assign _5136 = _1055 & _408;
    assign _5141 = _5136 ? _599 : _5140;
    assign _353 = _5141;
    always @(posedge _416) begin
        if (_414)
            _602 <= _5492;
        else
            _602 <= _353;
    end
    assign _3450 = { gnd,
                     _602 };
    assign _3452 = _3450 < _3451;
    assign _5143 = _3452 ? _602 : _599;
    assign _3449 = _1064[0:0];
    assign _5145 = _3449 ? _5144 : _5143;
    assign _5146 = _1058 ? _5145 : _599;
    assign _5142 = _1055 & _408;
    assign _5147 = _5142 ? _596 : _5146;
    assign _354 = _5147;
    always @(posedge _416) begin
        if (_414)
            _599 <= _5492;
        else
            _599 <= _354;
    end
    assign _3473 = { gnd,
                     _599 };
    assign _3475 = _3473 < _3474;
    assign _5150 = _3475 ? _599 : _596;
    assign _3467 = { gnd,
                     _593 };
    assign _3466 = { gnd,
                     _596 };
    assign _3468 = _3466 < _3467;
    assign _5149 = _3468 ? _593 : _596;
    assign _3465 = _1064[0:0];
    assign _5151 = _3465 ? _5150 : _5149;
    assign _5152 = _1058 ? _5151 : _596;
    assign _5148 = _1055 & _408;
    assign _5153 = _5148 ? _593 : _5152;
    assign _355 = _5153;
    always @(posedge _416) begin
        if (_414)
            _596 <= _5492;
        else
            _596 <= _355;
    end
    assign _3482 = { gnd,
                     _596 };
    assign _3484 = _3482 < _3483;
    assign _5155 = _3484 ? _596 : _593;
    assign _3481 = _1064[0:0];
    assign _5157 = _3481 ? _5156 : _5155;
    assign _5158 = _1058 ? _5157 : _593;
    assign _5154 = _1055 & _408;
    assign _5159 = _5154 ? _590 : _5158;
    assign _356 = _5159;
    always @(posedge _416) begin
        if (_414)
            _593 <= _5492;
        else
            _593 <= _356;
    end
    assign _3505 = { gnd,
                     _593 };
    assign _3507 = _3505 < _3506;
    assign _5162 = _3507 ? _593 : _590;
    assign _3499 = { gnd,
                     _587 };
    assign _3498 = { gnd,
                     _590 };
    assign _3500 = _3498 < _3499;
    assign _5161 = _3500 ? _587 : _590;
    assign _3497 = _1064[0:0];
    assign _5163 = _3497 ? _5162 : _5161;
    assign _5164 = _1058 ? _5163 : _590;
    assign _5160 = _1055 & _408;
    assign _5165 = _5160 ? _587 : _5164;
    assign _357 = _5165;
    always @(posedge _416) begin
        if (_414)
            _590 <= _5492;
        else
            _590 <= _357;
    end
    assign _3514 = { gnd,
                     _590 };
    assign _3516 = _3514 < _3515;
    assign _5167 = _3516 ? _590 : _587;
    assign _3513 = _1064[0:0];
    assign _5169 = _3513 ? _5168 : _5167;
    assign _5170 = _1058 ? _5169 : _587;
    assign _5166 = _1055 & _408;
    assign _5171 = _5166 ? _584 : _5170;
    assign _358 = _5171;
    always @(posedge _416) begin
        if (_414)
            _587 <= _5492;
        else
            _587 <= _358;
    end
    assign _3537 = { gnd,
                     _587 };
    assign _3539 = _3537 < _3538;
    assign _5174 = _3539 ? _587 : _584;
    assign _3531 = { gnd,
                     _581 };
    assign _3530 = { gnd,
                     _584 };
    assign _3532 = _3530 < _3531;
    assign _5173 = _3532 ? _581 : _584;
    assign _3529 = _1064[0:0];
    assign _5175 = _3529 ? _5174 : _5173;
    assign _5176 = _1058 ? _5175 : _584;
    assign _5172 = _1055 & _408;
    assign _5177 = _5172 ? _581 : _5176;
    assign _359 = _5177;
    always @(posedge _416) begin
        if (_414)
            _584 <= _5492;
        else
            _584 <= _359;
    end
    assign _3546 = { gnd,
                     _584 };
    assign _3548 = _3546 < _3547;
    assign _5179 = _3548 ? _584 : _581;
    assign _3545 = _1064[0:0];
    assign _5181 = _3545 ? _5180 : _5179;
    assign _5182 = _1058 ? _5181 : _581;
    assign _5178 = _1055 & _408;
    assign _5183 = _5178 ? _578 : _5182;
    assign _360 = _5183;
    always @(posedge _416) begin
        if (_414)
            _581 <= _5492;
        else
            _581 <= _360;
    end
    assign _3569 = { gnd,
                     _581 };
    assign _3571 = _3569 < _3570;
    assign _5186 = _3571 ? _581 : _578;
    assign _3563 = { gnd,
                     _575 };
    assign _3562 = { gnd,
                     _578 };
    assign _3564 = _3562 < _3563;
    assign _5185 = _3564 ? _575 : _578;
    assign _3561 = _1064[0:0];
    assign _5187 = _3561 ? _5186 : _5185;
    assign _5188 = _1058 ? _5187 : _578;
    assign _5184 = _1055 & _408;
    assign _5189 = _5184 ? _575 : _5188;
    assign _361 = _5189;
    always @(posedge _416) begin
        if (_414)
            _578 <= _5492;
        else
            _578 <= _361;
    end
    assign _3578 = { gnd,
                     _578 };
    assign _3580 = _3578 < _3579;
    assign _5191 = _3580 ? _578 : _575;
    assign _3577 = _1064[0:0];
    assign _5193 = _3577 ? _5192 : _5191;
    assign _5194 = _1058 ? _5193 : _575;
    assign _5190 = _1055 & _408;
    assign _5195 = _5190 ? _572 : _5194;
    assign _362 = _5195;
    always @(posedge _416) begin
        if (_414)
            _575 <= _5492;
        else
            _575 <= _362;
    end
    assign _3601 = { gnd,
                     _575 };
    assign _3603 = _3601 < _3602;
    assign _5198 = _3603 ? _575 : _572;
    assign _3595 = { gnd,
                     _569 };
    assign _3594 = { gnd,
                     _572 };
    assign _3596 = _3594 < _3595;
    assign _5197 = _3596 ? _569 : _572;
    assign _3593 = _1064[0:0];
    assign _5199 = _3593 ? _5198 : _5197;
    assign _5200 = _1058 ? _5199 : _572;
    assign _5196 = _1055 & _408;
    assign _5201 = _5196 ? _569 : _5200;
    assign _363 = _5201;
    always @(posedge _416) begin
        if (_414)
            _572 <= _5492;
        else
            _572 <= _363;
    end
    assign _3610 = { gnd,
                     _572 };
    assign _3612 = _3610 < _3611;
    assign _5203 = _3612 ? _572 : _569;
    assign _3609 = _1064[0:0];
    assign _5205 = _3609 ? _5204 : _5203;
    assign _5206 = _1058 ? _5205 : _569;
    assign _5202 = _1055 & _408;
    assign _5207 = _5202 ? _566 : _5206;
    assign _364 = _5207;
    always @(posedge _416) begin
        if (_414)
            _569 <= _5492;
        else
            _569 <= _364;
    end
    assign _3633 = { gnd,
                     _569 };
    assign _3635 = _3633 < _3634;
    assign _5210 = _3635 ? _569 : _566;
    assign _3627 = { gnd,
                     _563 };
    assign _3626 = { gnd,
                     _566 };
    assign _3628 = _3626 < _3627;
    assign _5209 = _3628 ? _563 : _566;
    assign _3625 = _1064[0:0];
    assign _5211 = _3625 ? _5210 : _5209;
    assign _5212 = _1058 ? _5211 : _566;
    assign _5208 = _1055 & _408;
    assign _5213 = _5208 ? _563 : _5212;
    assign _365 = _5213;
    always @(posedge _416) begin
        if (_414)
            _566 <= _5492;
        else
            _566 <= _365;
    end
    assign _3642 = { gnd,
                     _566 };
    assign _3644 = _3642 < _3643;
    assign _5215 = _3644 ? _566 : _563;
    assign _3641 = _1064[0:0];
    assign _5217 = _3641 ? _5216 : _5215;
    assign _5218 = _1058 ? _5217 : _563;
    assign _5214 = _1055 & _408;
    assign _5219 = _5214 ? _560 : _5218;
    assign _366 = _5219;
    always @(posedge _416) begin
        if (_414)
            _563 <= _5492;
        else
            _563 <= _366;
    end
    assign _3665 = { gnd,
                     _563 };
    assign _3667 = _3665 < _3666;
    assign _5222 = _3667 ? _563 : _560;
    assign _3659 = { gnd,
                     _557 };
    assign _3658 = { gnd,
                     _560 };
    assign _3660 = _3658 < _3659;
    assign _5221 = _3660 ? _557 : _560;
    assign _3657 = _1064[0:0];
    assign _5223 = _3657 ? _5222 : _5221;
    assign _5224 = _1058 ? _5223 : _560;
    assign _5220 = _1055 & _408;
    assign _5225 = _5220 ? _557 : _5224;
    assign _367 = _5225;
    always @(posedge _416) begin
        if (_414)
            _560 <= _5492;
        else
            _560 <= _367;
    end
    assign _3674 = { gnd,
                     _560 };
    assign _3676 = _3674 < _3675;
    assign _5227 = _3676 ? _560 : _557;
    assign _3673 = _1064[0:0];
    assign _5229 = _3673 ? _5228 : _5227;
    assign _5230 = _1058 ? _5229 : _557;
    assign _5226 = _1055 & _408;
    assign _5231 = _5226 ? _554 : _5230;
    assign _368 = _5231;
    always @(posedge _416) begin
        if (_414)
            _557 <= _5492;
        else
            _557 <= _368;
    end
    assign _3697 = { gnd,
                     _557 };
    assign _3699 = _3697 < _3698;
    assign _5234 = _3699 ? _557 : _554;
    assign _3691 = { gnd,
                     _551 };
    assign _3690 = { gnd,
                     _554 };
    assign _3692 = _3690 < _3691;
    assign _5233 = _3692 ? _551 : _554;
    assign _3689 = _1064[0:0];
    assign _5235 = _3689 ? _5234 : _5233;
    assign _5236 = _1058 ? _5235 : _554;
    assign _5232 = _1055 & _408;
    assign _5237 = _5232 ? _551 : _5236;
    assign _369 = _5237;
    always @(posedge _416) begin
        if (_414)
            _554 <= _5492;
        else
            _554 <= _369;
    end
    assign _3706 = { gnd,
                     _554 };
    assign _3708 = _3706 < _3707;
    assign _5239 = _3708 ? _554 : _551;
    assign _3705 = _1064[0:0];
    assign _5241 = _3705 ? _5240 : _5239;
    assign _5242 = _1058 ? _5241 : _551;
    assign _5238 = _1055 & _408;
    assign _5243 = _5238 ? _548 : _5242;
    assign _370 = _5243;
    always @(posedge _416) begin
        if (_414)
            _551 <= _5492;
        else
            _551 <= _370;
    end
    assign _3729 = { gnd,
                     _551 };
    assign _3731 = _3729 < _3730;
    assign _5246 = _3731 ? _551 : _548;
    assign _3723 = { gnd,
                     _545 };
    assign _3722 = { gnd,
                     _548 };
    assign _3724 = _3722 < _3723;
    assign _5245 = _3724 ? _545 : _548;
    assign _3721 = _1064[0:0];
    assign _5247 = _3721 ? _5246 : _5245;
    assign _5248 = _1058 ? _5247 : _548;
    assign _5244 = _1055 & _408;
    assign _5249 = _5244 ? _545 : _5248;
    assign _371 = _5249;
    always @(posedge _416) begin
        if (_414)
            _548 <= _5492;
        else
            _548 <= _371;
    end
    assign _3738 = { gnd,
                     _548 };
    assign _3740 = _3738 < _3739;
    assign _5251 = _3740 ? _548 : _545;
    assign _3737 = _1064[0:0];
    assign _5253 = _3737 ? _5252 : _5251;
    assign _5254 = _1058 ? _5253 : _545;
    assign _5250 = _1055 & _408;
    assign _5255 = _5250 ? _542 : _5254;
    assign _372 = _5255;
    always @(posedge _416) begin
        if (_414)
            _545 <= _5492;
        else
            _545 <= _372;
    end
    assign _3761 = { gnd,
                     _545 };
    assign _3763 = _3761 < _3762;
    assign _5258 = _3763 ? _545 : _542;
    assign _3755 = { gnd,
                     _539 };
    assign _3754 = { gnd,
                     _542 };
    assign _3756 = _3754 < _3755;
    assign _5257 = _3756 ? _539 : _542;
    assign _3753 = _1064[0:0];
    assign _5259 = _3753 ? _5258 : _5257;
    assign _5260 = _1058 ? _5259 : _542;
    assign _5256 = _1055 & _408;
    assign _5261 = _5256 ? _539 : _5260;
    assign _373 = _5261;
    always @(posedge _416) begin
        if (_414)
            _542 <= _5492;
        else
            _542 <= _373;
    end
    assign _3770 = { gnd,
                     _542 };
    assign _3772 = _3770 < _3771;
    assign _5263 = _3772 ? _542 : _539;
    assign _3769 = _1064[0:0];
    assign _5265 = _3769 ? _5264 : _5263;
    assign _5266 = _1058 ? _5265 : _539;
    assign _5262 = _1055 & _408;
    assign _5267 = _5262 ? _536 : _5266;
    assign _374 = _5267;
    always @(posedge _416) begin
        if (_414)
            _539 <= _5492;
        else
            _539 <= _374;
    end
    assign _3793 = { gnd,
                     _539 };
    assign _3795 = _3793 < _3794;
    assign _5270 = _3795 ? _539 : _536;
    assign _3787 = { gnd,
                     _533 };
    assign _3786 = { gnd,
                     _536 };
    assign _3788 = _3786 < _3787;
    assign _5269 = _3788 ? _533 : _536;
    assign _3785 = _1064[0:0];
    assign _5271 = _3785 ? _5270 : _5269;
    assign _5272 = _1058 ? _5271 : _536;
    assign _5268 = _1055 & _408;
    assign _5273 = _5268 ? _533 : _5272;
    assign _375 = _5273;
    always @(posedge _416) begin
        if (_414)
            _536 <= _5492;
        else
            _536 <= _375;
    end
    assign _3802 = { gnd,
                     _536 };
    assign _3804 = _3802 < _3803;
    assign _5275 = _3804 ? _536 : _533;
    assign _3801 = _1064[0:0];
    assign _5277 = _3801 ? _5276 : _5275;
    assign _5278 = _1058 ? _5277 : _533;
    assign _5274 = _1055 & _408;
    assign _5279 = _5274 ? _530 : _5278;
    assign _376 = _5279;
    always @(posedge _416) begin
        if (_414)
            _533 <= _5492;
        else
            _533 <= _376;
    end
    assign _3825 = { gnd,
                     _533 };
    assign _3827 = _3825 < _3826;
    assign _5282 = _3827 ? _533 : _530;
    assign _3819 = { gnd,
                     _527 };
    assign _3818 = { gnd,
                     _530 };
    assign _3820 = _3818 < _3819;
    assign _5281 = _3820 ? _527 : _530;
    assign _3817 = _1064[0:0];
    assign _5283 = _3817 ? _5282 : _5281;
    assign _5284 = _1058 ? _5283 : _530;
    assign _5280 = _1055 & _408;
    assign _5285 = _5280 ? _527 : _5284;
    assign _377 = _5285;
    always @(posedge _416) begin
        if (_414)
            _530 <= _5492;
        else
            _530 <= _377;
    end
    assign _3834 = { gnd,
                     _530 };
    assign _3836 = _3834 < _3835;
    assign _5287 = _3836 ? _530 : _527;
    assign _3833 = _1064[0:0];
    assign _5289 = _3833 ? _5288 : _5287;
    assign _5290 = _1058 ? _5289 : _527;
    assign _5286 = _1055 & _408;
    assign _5291 = _5286 ? _524 : _5290;
    assign _378 = _5291;
    always @(posedge _416) begin
        if (_414)
            _527 <= _5492;
        else
            _527 <= _378;
    end
    assign _3857 = { gnd,
                     _527 };
    assign _3859 = _3857 < _3858;
    assign _5294 = _3859 ? _527 : _524;
    assign _3851 = { gnd,
                     _521 };
    assign _3850 = { gnd,
                     _524 };
    assign _3852 = _3850 < _3851;
    assign _5293 = _3852 ? _521 : _524;
    assign _3849 = _1064[0:0];
    assign _5295 = _3849 ? _5294 : _5293;
    assign _5296 = _1058 ? _5295 : _524;
    assign _5292 = _1055 & _408;
    assign _5297 = _5292 ? _521 : _5296;
    assign _379 = _5297;
    always @(posedge _416) begin
        if (_414)
            _524 <= _5492;
        else
            _524 <= _379;
    end
    assign _3866 = { gnd,
                     _524 };
    assign _3868 = _3866 < _3867;
    assign _5299 = _3868 ? _524 : _521;
    assign _3865 = _1064[0:0];
    assign _5301 = _3865 ? _5300 : _5299;
    assign _5302 = _1058 ? _5301 : _521;
    assign _5298 = _1055 & _408;
    assign _5303 = _5298 ? _518 : _5302;
    assign _380 = _5303;
    always @(posedge _416) begin
        if (_414)
            _521 <= _5492;
        else
            _521 <= _380;
    end
    assign _3889 = { gnd,
                     _521 };
    assign _3891 = _3889 < _3890;
    assign _5306 = _3891 ? _521 : _518;
    assign _3883 = { gnd,
                     _515 };
    assign _3882 = { gnd,
                     _518 };
    assign _3884 = _3882 < _3883;
    assign _5305 = _3884 ? _515 : _518;
    assign _3881 = _1064[0:0];
    assign _5307 = _3881 ? _5306 : _5305;
    assign _5308 = _1058 ? _5307 : _518;
    assign _5304 = _1055 & _408;
    assign _5309 = _5304 ? _515 : _5308;
    assign _381 = _5309;
    always @(posedge _416) begin
        if (_414)
            _518 <= _5492;
        else
            _518 <= _381;
    end
    assign _3898 = { gnd,
                     _518 };
    assign _3900 = _3898 < _3899;
    assign _5311 = _3900 ? _518 : _515;
    assign _3897 = _1064[0:0];
    assign _5313 = _3897 ? _5312 : _5311;
    assign _5314 = _1058 ? _5313 : _515;
    assign _5310 = _1055 & _408;
    assign _5315 = _5310 ? _512 : _5314;
    assign _382 = _5315;
    always @(posedge _416) begin
        if (_414)
            _515 <= _5492;
        else
            _515 <= _382;
    end
    assign _3921 = { gnd,
                     _515 };
    assign _3923 = _3921 < _3922;
    assign _5318 = _3923 ? _515 : _512;
    assign _3915 = { gnd,
                     _509 };
    assign _3914 = { gnd,
                     _512 };
    assign _3916 = _3914 < _3915;
    assign _5317 = _3916 ? _509 : _512;
    assign _3913 = _1064[0:0];
    assign _5319 = _3913 ? _5318 : _5317;
    assign _5320 = _1058 ? _5319 : _512;
    assign _5316 = _1055 & _408;
    assign _5321 = _5316 ? _509 : _5320;
    assign _383 = _5321;
    always @(posedge _416) begin
        if (_414)
            _512 <= _5492;
        else
            _512 <= _383;
    end
    assign _3930 = { gnd,
                     _512 };
    assign _3932 = _3930 < _3931;
    assign _5323 = _3932 ? _512 : _509;
    assign _3929 = _1064[0:0];
    assign _5325 = _3929 ? _5324 : _5323;
    assign _5326 = _1058 ? _5325 : _509;
    assign _5322 = _1055 & _408;
    assign _5327 = _5322 ? _506 : _5326;
    assign _384 = _5327;
    always @(posedge _416) begin
        if (_414)
            _509 <= _5492;
        else
            _509 <= _384;
    end
    assign _3953 = { gnd,
                     _509 };
    assign _3955 = _3953 < _3954;
    assign _5330 = _3955 ? _509 : _506;
    assign _3947 = { gnd,
                     _503 };
    assign _3946 = { gnd,
                     _506 };
    assign _3948 = _3946 < _3947;
    assign _5329 = _3948 ? _503 : _506;
    assign _3945 = _1064[0:0];
    assign _5331 = _3945 ? _5330 : _5329;
    assign _5332 = _1058 ? _5331 : _506;
    assign _5328 = _1055 & _408;
    assign _5333 = _5328 ? _503 : _5332;
    assign _385 = _5333;
    always @(posedge _416) begin
        if (_414)
            _506 <= _5492;
        else
            _506 <= _385;
    end
    assign _3962 = { gnd,
                     _506 };
    assign _3964 = _3962 < _3963;
    assign _5335 = _3964 ? _506 : _503;
    assign _3961 = _1064[0:0];
    assign _5337 = _3961 ? _5336 : _5335;
    assign _5338 = _1058 ? _5337 : _503;
    assign _5334 = _1055 & _408;
    assign _5339 = _5334 ? _500 : _5338;
    assign _386 = _5339;
    always @(posedge _416) begin
        if (_414)
            _503 <= _5492;
        else
            _503 <= _386;
    end
    assign _3985 = { gnd,
                     _503 };
    assign _3987 = _3985 < _3986;
    assign _5342 = _3987 ? _503 : _500;
    assign _3979 = { gnd,
                     _497 };
    assign _3978 = { gnd,
                     _500 };
    assign _3980 = _3978 < _3979;
    assign _5341 = _3980 ? _497 : _500;
    assign _3977 = _1064[0:0];
    assign _5343 = _3977 ? _5342 : _5341;
    assign _5344 = _1058 ? _5343 : _500;
    assign _5340 = _1055 & _408;
    assign _5345 = _5340 ? _497 : _5344;
    assign _387 = _5345;
    always @(posedge _416) begin
        if (_414)
            _500 <= _5492;
        else
            _500 <= _387;
    end
    assign _3994 = { gnd,
                     _500 };
    assign _3996 = _3994 < _3995;
    assign _5347 = _3996 ? _500 : _497;
    assign _3993 = _1064[0:0];
    assign _5349 = _3993 ? _5348 : _5347;
    assign _5350 = _1058 ? _5349 : _497;
    assign _5346 = _1055 & _408;
    assign _5351 = _5346 ? _494 : _5350;
    assign _388 = _5351;
    always @(posedge _416) begin
        if (_414)
            _497 <= _5492;
        else
            _497 <= _388;
    end
    assign _4017 = { gnd,
                     _497 };
    assign _4019 = _4017 < _4018;
    assign _5354 = _4019 ? _497 : _494;
    assign _4011 = { gnd,
                     _491 };
    assign _4010 = { gnd,
                     _494 };
    assign _4012 = _4010 < _4011;
    assign _5353 = _4012 ? _491 : _494;
    assign _4009 = _1064[0:0];
    assign _5355 = _4009 ? _5354 : _5353;
    assign _5356 = _1058 ? _5355 : _494;
    assign _5352 = _1055 & _408;
    assign _5357 = _5352 ? _491 : _5356;
    assign _389 = _5357;
    always @(posedge _416) begin
        if (_414)
            _494 <= _5492;
        else
            _494 <= _389;
    end
    assign _4026 = { gnd,
                     _494 };
    assign _4028 = _4026 < _4027;
    assign _5359 = _4028 ? _494 : _491;
    assign _4025 = _1064[0:0];
    assign _5361 = _4025 ? _5360 : _5359;
    assign _5362 = _1058 ? _5361 : _491;
    assign _5358 = _1055 & _408;
    assign _5363 = _5358 ? _488 : _5362;
    assign _390 = _5363;
    always @(posedge _416) begin
        if (_414)
            _491 <= _5492;
        else
            _491 <= _390;
    end
    assign _4049 = { gnd,
                     _491 };
    assign _4051 = _4049 < _4050;
    assign _5366 = _4051 ? _491 : _488;
    assign _4043 = { gnd,
                     _485 };
    assign _4042 = { gnd,
                     _488 };
    assign _4044 = _4042 < _4043;
    assign _5365 = _4044 ? _485 : _488;
    assign _4041 = _1064[0:0];
    assign _5367 = _4041 ? _5366 : _5365;
    assign _5368 = _1058 ? _5367 : _488;
    assign _5364 = _1055 & _408;
    assign _5369 = _5364 ? _485 : _5368;
    assign _391 = _5369;
    always @(posedge _416) begin
        if (_414)
            _488 <= _5492;
        else
            _488 <= _391;
    end
    assign _4058 = { gnd,
                     _488 };
    assign _4060 = _4058 < _4059;
    assign _5371 = _4060 ? _488 : _485;
    assign _4057 = _1064[0:0];
    assign _5373 = _4057 ? _5372 : _5371;
    assign _5374 = _1058 ? _5373 : _485;
    assign _5370 = _1055 & _408;
    assign _5375 = _5370 ? _482 : _5374;
    assign _392 = _5375;
    always @(posedge _416) begin
        if (_414)
            _485 <= _5492;
        else
            _485 <= _392;
    end
    assign _4081 = { gnd,
                     _485 };
    assign _4083 = _4081 < _4082;
    assign _5378 = _4083 ? _485 : _482;
    assign _4075 = { gnd,
                     _479 };
    assign _4074 = { gnd,
                     _482 };
    assign _4076 = _4074 < _4075;
    assign _5377 = _4076 ? _479 : _482;
    assign _4073 = _1064[0:0];
    assign _5379 = _4073 ? _5378 : _5377;
    assign _5380 = _1058 ? _5379 : _482;
    assign _5376 = _1055 & _408;
    assign _5381 = _5376 ? _479 : _5380;
    assign _393 = _5381;
    always @(posedge _416) begin
        if (_414)
            _482 <= _5492;
        else
            _482 <= _393;
    end
    assign _4090 = { gnd,
                     _482 };
    assign _4092 = _4090 < _4091;
    assign _5383 = _4092 ? _482 : _479;
    assign _4089 = _1064[0:0];
    assign _5385 = _4089 ? _5384 : _5383;
    assign _5386 = _1058 ? _5385 : _479;
    assign _5382 = _1055 & _408;
    assign _5387 = _5382 ? _476 : _5386;
    assign _394 = _5387;
    always @(posedge _416) begin
        if (_414)
            _479 <= _5492;
        else
            _479 <= _394;
    end
    assign _4113 = { gnd,
                     _479 };
    assign _4115 = _4113 < _4114;
    assign _5390 = _4115 ? _479 : _476;
    assign _4107 = { gnd,
                     _473 };
    assign _4106 = { gnd,
                     _476 };
    assign _4108 = _4106 < _4107;
    assign _5389 = _4108 ? _473 : _476;
    assign _4105 = _1064[0:0];
    assign _5391 = _4105 ? _5390 : _5389;
    assign _5392 = _1058 ? _5391 : _476;
    assign _5388 = _1055 & _408;
    assign _5393 = _5388 ? _473 : _5392;
    assign _395 = _5393;
    always @(posedge _416) begin
        if (_414)
            _476 <= _5492;
        else
            _476 <= _395;
    end
    assign _4122 = { gnd,
                     _476 };
    assign _4124 = _4122 < _4123;
    assign _5395 = _4124 ? _476 : _473;
    assign _4121 = _1064[0:0];
    assign _5397 = _4121 ? _5396 : _5395;
    assign _5398 = _1058 ? _5397 : _473;
    assign _5394 = _1055 & _408;
    assign _5399 = _5394 ? _470 : _5398;
    assign _396 = _5399;
    always @(posedge _416) begin
        if (_414)
            _473 <= _5492;
        else
            _473 <= _396;
    end
    assign _4145 = { gnd,
                     _473 };
    assign _4147 = _4145 < _4146;
    assign _5402 = _4147 ? _473 : _470;
    assign _4139 = { gnd,
                     _467 };
    assign _4138 = { gnd,
                     _470 };
    assign _4140 = _4138 < _4139;
    assign _5401 = _4140 ? _467 : _470;
    assign _4137 = _1064[0:0];
    assign _5403 = _4137 ? _5402 : _5401;
    assign _5404 = _1058 ? _5403 : _470;
    assign _5400 = _1055 & _408;
    assign _5405 = _5400 ? _467 : _5404;
    assign _397 = _5405;
    always @(posedge _416) begin
        if (_414)
            _470 <= _5492;
        else
            _470 <= _397;
    end
    assign _4154 = { gnd,
                     _470 };
    assign _4156 = _4154 < _4155;
    assign _5407 = _4156 ? _470 : _467;
    assign _4153 = _1064[0:0];
    assign _5409 = _4153 ? _5408 : _5407;
    assign _5410 = _1058 ? _5409 : _467;
    assign _5406 = _1055 & _408;
    assign _5411 = _5406 ? _464 : _5410;
    assign _398 = _5411;
    always @(posedge _416) begin
        if (_414)
            _467 <= _5492;
        else
            _467 <= _398;
    end
    assign _4177 = { gnd,
                     _467 };
    assign _4179 = _4177 < _4178;
    assign _5414 = _4179 ? _467 : _464;
    assign _4171 = { gnd,
                     _461 };
    assign _4170 = { gnd,
                     _464 };
    assign _4172 = _4170 < _4171;
    assign _5413 = _4172 ? _461 : _464;
    assign _4169 = _1064[0:0];
    assign _5415 = _4169 ? _5414 : _5413;
    assign _5416 = _1058 ? _5415 : _464;
    assign _5412 = _1055 & _408;
    assign _5417 = _5412 ? _461 : _5416;
    assign _399 = _5417;
    always @(posedge _416) begin
        if (_414)
            _464 <= _5492;
        else
            _464 <= _399;
    end
    assign _4186 = { gnd,
                     _464 };
    assign _4188 = _4186 < _4187;
    assign _5419 = _4188 ? _464 : _461;
    assign _4185 = _1064[0:0];
    assign _5421 = _4185 ? _5420 : _5419;
    assign _5422 = _1058 ? _5421 : _461;
    assign _5418 = _1055 & _408;
    assign _5423 = _5418 ? _458 : _5422;
    assign _400 = _5423;
    always @(posedge _416) begin
        if (_414)
            _461 <= _5492;
        else
            _461 <= _400;
    end
    assign _4209 = { gnd,
                     _461 };
    assign _4211 = _4209 < _4210;
    assign _5426 = _4211 ? _461 : _458;
    assign _4203 = { gnd,
                     _455 };
    assign _4202 = { gnd,
                     _458 };
    assign _4204 = _4202 < _4203;
    assign _5425 = _4204 ? _455 : _458;
    assign _4201 = _1064[0:0];
    assign _5427 = _4201 ? _5426 : _5425;
    assign _5428 = _1058 ? _5427 : _458;
    assign _5424 = _1055 & _408;
    assign _5429 = _5424 ? _455 : _5428;
    assign _401 = _5429;
    always @(posedge _416) begin
        if (_414)
            _458 <= _5492;
        else
            _458 <= _401;
    end
    assign _4218 = { gnd,
                     _458 };
    assign _4220 = _4218 < _4219;
    assign _5431 = _4220 ? _458 : _455;
    assign _4217 = _1064[0:0];
    assign _5433 = _4217 ? _5432 : _5431;
    assign _5434 = _1058 ? _5433 : _455;
    assign _5430 = _1055 & _408;
    assign _5435 = _5430 ? _452 : _5434;
    assign _402 = _5435;
    always @(posedge _416) begin
        if (_414)
            _455 <= _5492;
        else
            _455 <= _402;
    end
    assign _4241 = { gnd,
                     _455 };
    assign _4243 = _4241 < _4242;
    assign _5451 = _4243 ? _455 : _452;
    assign _404 = wr_start;
    assign _5443 = { gnd,
                     _449 };
    assign _5442 = { gnd,
                     _449 };
    assign _5444 = _5442 < _5443;
    assign _5445 = _5444 ? _449 : _449;
    assign _5441 = _5440 ? _452 : _449;
    assign _5446 = _5437 ? _5445 : _5441;
    assign _5447 = _1058 ? _5446 : _449;
    assign _5436 = _1055 & _408;
    assign _5448 = _5436 ? _404 : _5447;
    assign _405 = _5448;
    always @(posedge _416) begin
        if (_414)
            _449 <= _5492;
        else
            _449 <= _405;
    end
    assign _4235 = { gnd,
                     _449 };
    assign _4234 = { gnd,
                     _452 };
    assign _4236 = _4234 < _4235;
    assign _5450 = _4236 ? _449 : _452;
    assign _4233 = _1064[0:0];
    assign _5452 = _4233 ? _5451 : _5450;
    assign _5453 = _1058 ? _5452 : _452;
    assign _5449 = _1055 & _408;
    assign _5454 = _5449 ? _449 : _5453;
    assign _406 = _5454;
    always @(posedge _416) begin
        if (_414)
            _452 <= _5492;
        else
            _452 <= _406;
    end
    assign _5438 = { gnd,
                     _452 };
    assign _5440 = _5438 < _5439;
    assign _5456 = _5440 ? _4227 : _4239;
    assign _5437 = _1064[0:0];
    assign _5458 = _5437 ? _5457 : _5456;
    assign _5459 = _1058 ? _5458 : _4239;
    assign _408 = wr_enable;
    assign _1055 = _426 == _424;
    assign _5455 = _1055 & _408;
    assign _5460 = _5455 ? _5 : _5459;
    assign _409 = _5460;
    always @(posedge _416) begin
        if (_414)
            _4239 <= _5492;
        else
            _4239 <= _409;
    end
    always @* begin
        case (_446)
        0:
            _5462 <= _4239;
        1:
            _5462 <= _4227;
        2:
            _5462 <= _4207;
        3:
            _5462 <= _4195;
        4:
            _5462 <= _4175;
        5:
            _5462 <= _4163;
        6:
            _5462 <= _4143;
        7:
            _5462 <= _4131;
        8:
            _5462 <= _4111;
        9:
            _5462 <= _4099;
        10:
            _5462 <= _4079;
        11:
            _5462 <= _4067;
        12:
            _5462 <= _4047;
        13:
            _5462 <= _4035;
        14:
            _5462 <= _4015;
        15:
            _5462 <= _4003;
        16:
            _5462 <= _3983;
        17:
            _5462 <= _3971;
        18:
            _5462 <= _3951;
        19:
            _5462 <= _3939;
        20:
            _5462 <= _3919;
        21:
            _5462 <= _3907;
        22:
            _5462 <= _3887;
        23:
            _5462 <= _3875;
        24:
            _5462 <= _3855;
        25:
            _5462 <= _3843;
        26:
            _5462 <= _3823;
        27:
            _5462 <= _3811;
        28:
            _5462 <= _3791;
        29:
            _5462 <= _3779;
        30:
            _5462 <= _3759;
        31:
            _5462 <= _3747;
        32:
            _5462 <= _3727;
        33:
            _5462 <= _3715;
        34:
            _5462 <= _3695;
        35:
            _5462 <= _3683;
        36:
            _5462 <= _3663;
        37:
            _5462 <= _3651;
        38:
            _5462 <= _3631;
        39:
            _5462 <= _3619;
        40:
            _5462 <= _3599;
        41:
            _5462 <= _3587;
        42:
            _5462 <= _3567;
        43:
            _5462 <= _3555;
        44:
            _5462 <= _3535;
        45:
            _5462 <= _3523;
        46:
            _5462 <= _3503;
        47:
            _5462 <= _3491;
        48:
            _5462 <= _3471;
        49:
            _5462 <= _3459;
        50:
            _5462 <= _3439;
        51:
            _5462 <= _3427;
        52:
            _5462 <= _3407;
        53:
            _5462 <= _3395;
        54:
            _5462 <= _3375;
        55:
            _5462 <= _3363;
        56:
            _5462 <= _3343;
        57:
            _5462 <= _3331;
        58:
            _5462 <= _3311;
        59:
            _5462 <= _3299;
        60:
            _5462 <= _3279;
        61:
            _5462 <= _3267;
        62:
            _5462 <= _3247;
        63:
            _5462 <= _3235;
        64:
            _5462 <= _3215;
        65:
            _5462 <= _3203;
        66:
            _5462 <= _3183;
        67:
            _5462 <= _3171;
        68:
            _5462 <= _3151;
        69:
            _5462 <= _3139;
        70:
            _5462 <= _3119;
        71:
            _5462 <= _3107;
        72:
            _5462 <= _3087;
        73:
            _5462 <= _3075;
        74:
            _5462 <= _3055;
        75:
            _5462 <= _3043;
        76:
            _5462 <= _3023;
        77:
            _5462 <= _3011;
        78:
            _5462 <= _2991;
        79:
            _5462 <= _2979;
        80:
            _5462 <= _2959;
        81:
            _5462 <= _2947;
        82:
            _5462 <= _2927;
        83:
            _5462 <= _2915;
        84:
            _5462 <= _2895;
        85:
            _5462 <= _2883;
        86:
            _5462 <= _2863;
        87:
            _5462 <= _2851;
        88:
            _5462 <= _2831;
        89:
            _5462 <= _2819;
        90:
            _5462 <= _2799;
        91:
            _5462 <= _2787;
        92:
            _5462 <= _2767;
        93:
            _5462 <= _2755;
        94:
            _5462 <= _2735;
        95:
            _5462 <= _2723;
        96:
            _5462 <= _2703;
        97:
            _5462 <= _2691;
        98:
            _5462 <= _2671;
        99:
            _5462 <= _2659;
        100:
            _5462 <= _2639;
        101:
            _5462 <= _2627;
        102:
            _5462 <= _2607;
        103:
            _5462 <= _2595;
        104:
            _5462 <= _2575;
        105:
            _5462 <= _2563;
        106:
            _5462 <= _2543;
        107:
            _5462 <= _2531;
        108:
            _5462 <= _2511;
        109:
            _5462 <= _2499;
        110:
            _5462 <= _2479;
        111:
            _5462 <= _2467;
        112:
            _5462 <= _2447;
        113:
            _5462 <= _2435;
        114:
            _5462 <= _2415;
        115:
            _5462 <= _2403;
        116:
            _5462 <= _2383;
        117:
            _5462 <= _2371;
        118:
            _5462 <= _2351;
        119:
            _5462 <= _2339;
        120:
            _5462 <= _2319;
        121:
            _5462 <= _2307;
        122:
            _5462 <= _2287;
        123:
            _5462 <= _2275;
        124:
            _5462 <= _2255;
        125:
            _5462 <= _2243;
        126:
            _5462 <= _2223;
        127:
            _5462 <= _2211;
        128:
            _5462 <= _2191;
        129:
            _5462 <= _2179;
        130:
            _5462 <= _2159;
        131:
            _5462 <= _2147;
        132:
            _5462 <= _2127;
        133:
            _5462 <= _2115;
        134:
            _5462 <= _2095;
        135:
            _5462 <= _2083;
        136:
            _5462 <= _2063;
        137:
            _5462 <= _2051;
        138:
            _5462 <= _2031;
        139:
            _5462 <= _2019;
        140:
            _5462 <= _1999;
        141:
            _5462 <= _1987;
        142:
            _5462 <= _1967;
        143:
            _5462 <= _1955;
        144:
            _5462 <= _1935;
        145:
            _5462 <= _1923;
        146:
            _5462 <= _1903;
        147:
            _5462 <= _1891;
        148:
            _5462 <= _1871;
        149:
            _5462 <= _1859;
        150:
            _5462 <= _1839;
        151:
            _5462 <= _1827;
        152:
            _5462 <= _1807;
        153:
            _5462 <= _1795;
        154:
            _5462 <= _1775;
        155:
            _5462 <= _1763;
        156:
            _5462 <= _1743;
        157:
            _5462 <= _1731;
        158:
            _5462 <= _1711;
        159:
            _5462 <= _1699;
        160:
            _5462 <= _1679;
        161:
            _5462 <= _1667;
        162:
            _5462 <= _1647;
        163:
            _5462 <= _1635;
        164:
            _5462 <= _1615;
        165:
            _5462 <= _1603;
        166:
            _5462 <= _1583;
        167:
            _5462 <= _1571;
        168:
            _5462 <= _1551;
        169:
            _5462 <= _1539;
        170:
            _5462 <= _1519;
        171:
            _5462 <= _1507;
        172:
            _5462 <= _1487;
        173:
            _5462 <= _1475;
        174:
            _5462 <= _1455;
        175:
            _5462 <= _1443;
        176:
            _5462 <= _1423;
        177:
            _5462 <= _1411;
        178:
            _5462 <= _1391;
        179:
            _5462 <= _1379;
        180:
            _5462 <= _1359;
        181:
            _5462 <= _1347;
        182:
            _5462 <= _1327;
        183:
            _5462 <= _1315;
        184:
            _5462 <= _1295;
        185:
            _5462 <= _1283;
        186:
            _5462 <= _1263;
        187:
            _5462 <= _1251;
        188:
            _5462 <= _1231;
        189:
            _5462 <= _1219;
        190:
            _5462 <= _1199;
        191:
            _5462 <= _1187;
        192:
            _5462 <= _1167;
        193:
            _5462 <= _1155;
        194:
            _5462 <= _1135;
        195:
            _5462 <= _1123;
        196:
            _5462 <= _1103;
        197:
            _5462 <= _1091;
        198:
            _5462 <= _1071;
        default:
            _5462 <= _1061;
        endcase
    end
    assign _5461 = _436 & _1050;
    assign _5467 = _5461 ? _5466 : _5462;
    assign _5468 = _430 ? _5467 : _440;
    assign _410 = _5468;
    always @(posedge _416) begin
        if (_414)
            _440 <= _5492;
        else
            _440 <= _410;
    end
    assign _442 = _440 + _5495;
    assign _443 = { gnd,
                    _442 };
    assign _1049 = _443 < _1048;
    assign _1050 = ~ _1049;
    assign _5488 = ~ _1050;
    assign _5489 = _5488 | _5472;
    assign _435 = 1'b0;
    assign _5473 = _5472 ? gnd : _436;
    assign _5474 = _430 ? vdd : _5473;
    assign _411 = _5474;
    always @(posedge _416) begin
        if (_414)
            _436 <= _435;
        else
            _436 <= _411;
    end
    assign vdd = 1'b1;
    assign _424 = 2'b00;
    assign _427 = 2'b11;
    assign _5470 = 17'b00000000011001000;
    assign _445 = 16'b0000000000000000;
    assign _5475 = 16'b0000000000000001;
    assign _5476 = _446 + _5475;
    assign _412 = _5476;
    always @(posedge _416) begin
        if (_414)
            _446 <= _445;
        else
            if (_430)
                _446 <= _412;
    end
    assign _5469 = { gnd,
                     _446 };
    assign _5471 = _5469 < _5470;
    assign _5472 = ~ _5471;
    assign _5485 = _5472 ? _427 : _429;
    assign _429 = 2'b10;
    assign _1058 = _426 == _1057;
    assign _414 = clear;
    assign _416 = clock;
    assign _5478 = _1064 + _5475;
    assign _417 = _5478;
    always @(posedge _416) begin
        if (_414)
            _1064 <= _445;
        else
            if (_1058)
                _1064 <= _417;
    end
    assign gnd = 1'b0;
    assign _5480 = { gnd,
                     _1064 };
    assign _5482 = _5480 < _5470;
    assign _5483 = ~ _5482;
    assign _5484 = _5483 ? _429 : _1057;
    assign _1057 = 2'b01;
    assign _419 = start_processing;
    assign _5479 = _419 ? _1057 : _424;
    always @* begin
        case (_426)
        0:
            _5486 <= _5479;
        1:
            _5486 <= _5484;
        2:
            _5486 <= _5485;
        default:
            _5486 <= _427;
        endcase
    end
    assign _420 = _5486;
    always @(posedge _416) begin
        if (_414)
            _426 <= _424;
        else
            _426 <= _420;
    end
    assign _430 = _426 == _429;
    assign _5487 = _430 & _436;
    assign _5490 = _5487 & _5489;
    assign _5498 = _5490 ? _5497 : _5493;
    assign _421 = _5498;
    always @(posedge _416) begin
        if (_414)
            _5493 <= _5492;
        else
            _5493 <= _421;
    end
    assign result = _5493;
    assign done_flag = _428;
    assign state_debug = _426;

endmodule
